library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package multiple_access_ram_pkg is

    type addr_type is array (3 downto 0) of std_logic_vector(15 downto 0);
    type data_type is array (3 downto 0) of std_logic_vector(31 downto 0);

end package multiple_access_ram_pkg;

package body multiple_access_ram_pkg is

end package body multiple_access_ram_pkg;