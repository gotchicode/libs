library IEEE;                                                                 
use IEEE.std_logic_1164.all;                                                  
use IEEE.numeric_std.all;                                                     
                                                                              
entity test is                                                                  
 port (                                                                       
            clk             : in std_logic;                                   
            addr_in         : in std_logic_vector(7 downto 0);               
            rd_en           : in std_logic;                                   
                                                                              
            data_out        : out std_logic_vector(31 downto 0);              
            data_out_en     : out std_logic                                   
 );                                                                           
end entity test;                                                                
                                                                              
architecture rtl of test is                                                     
                                                                              
type ROM_type is array (0 to 255) of std_logic_vector(31 downto 0);            
signal ROM: ROM_type;                                                         
                                                                              
begin                                                                         
ROM(0) <= std_logic_vector(to_signed(0,32));
ROM(1) <= std_logic_vector(to_signed(25,32));
ROM(2) <= std_logic_vector(to_signed(50,32));
ROM(3) <= std_logic_vector(to_signed(75,32));
ROM(4) <= std_logic_vector(to_signed(100,32));
ROM(5) <= std_logic_vector(to_signed(125,32));
ROM(6) <= std_logic_vector(to_signed(150,32));
ROM(7) <= std_logic_vector(to_signed(175,32));
ROM(8) <= std_logic_vector(to_signed(200,32));
ROM(9) <= std_logic_vector(to_signed(224,32));
ROM(10) <= std_logic_vector(to_signed(249,32));
ROM(11) <= std_logic_vector(to_signed(273,32));
ROM(12) <= std_logic_vector(to_signed(297,32));
ROM(13) <= std_logic_vector(to_signed(321,32));
ROM(14) <= std_logic_vector(to_signed(345,32));
ROM(15) <= std_logic_vector(to_signed(369,32));
ROM(16) <= std_logic_vector(to_signed(392,32));
ROM(17) <= std_logic_vector(to_signed(415,32));
ROM(18) <= std_logic_vector(to_signed(438,32));
ROM(19) <= std_logic_vector(to_signed(460,32));
ROM(20) <= std_logic_vector(to_signed(483,32));
ROM(21) <= std_logic_vector(to_signed(505,32));
ROM(22) <= std_logic_vector(to_signed(526,32));
ROM(23) <= std_logic_vector(to_signed(548,32));
ROM(24) <= std_logic_vector(to_signed(569,32));
ROM(25) <= std_logic_vector(to_signed(590,32));
ROM(26) <= std_logic_vector(to_signed(610,32));
ROM(27) <= std_logic_vector(to_signed(630,32));
ROM(28) <= std_logic_vector(to_signed(650,32));
ROM(29) <= std_logic_vector(to_signed(669,32));
ROM(30) <= std_logic_vector(to_signed(688,32));
ROM(31) <= std_logic_vector(to_signed(706,32));
ROM(32) <= std_logic_vector(to_signed(724,32));
ROM(33) <= std_logic_vector(to_signed(742,32));
ROM(34) <= std_logic_vector(to_signed(759,32));
ROM(35) <= std_logic_vector(to_signed(775,32));
ROM(36) <= std_logic_vector(to_signed(792,32));
ROM(37) <= std_logic_vector(to_signed(807,32));
ROM(38) <= std_logic_vector(to_signed(822,32));
ROM(39) <= std_logic_vector(to_signed(837,32));
ROM(40) <= std_logic_vector(to_signed(851,32));
ROM(41) <= std_logic_vector(to_signed(865,32));
ROM(42) <= std_logic_vector(to_signed(878,32));
ROM(43) <= std_logic_vector(to_signed(891,32));
ROM(44) <= std_logic_vector(to_signed(903,32));
ROM(45) <= std_logic_vector(to_signed(915,32));
ROM(46) <= std_logic_vector(to_signed(926,32));
ROM(47) <= std_logic_vector(to_signed(936,32));
ROM(48) <= std_logic_vector(to_signed(946,32));
ROM(49) <= std_logic_vector(to_signed(955,32));
ROM(50) <= std_logic_vector(to_signed(964,32));
ROM(51) <= std_logic_vector(to_signed(972,32));
ROM(52) <= std_logic_vector(to_signed(980,32));
ROM(53) <= std_logic_vector(to_signed(987,32));
ROM(54) <= std_logic_vector(to_signed(993,32));
ROM(55) <= std_logic_vector(to_signed(999,32));
ROM(56) <= std_logic_vector(to_signed(1004,32));
ROM(57) <= std_logic_vector(to_signed(1009,32));
ROM(58) <= std_logic_vector(to_signed(1013,32));
ROM(59) <= std_logic_vector(to_signed(1016,32));
ROM(60) <= std_logic_vector(to_signed(1019,32));
ROM(61) <= std_logic_vector(to_signed(1021,32));
ROM(62) <= std_logic_vector(to_signed(1023,32));
ROM(63) <= std_logic_vector(to_signed(1024,32));
ROM(64) <= std_logic_vector(to_signed(1024,32));
ROM(65) <= std_logic_vector(to_signed(1024,32));
ROM(66) <= std_logic_vector(to_signed(1023,32));
ROM(67) <= std_logic_vector(to_signed(1021,32));
ROM(68) <= std_logic_vector(to_signed(1019,32));
ROM(69) <= std_logic_vector(to_signed(1016,32));
ROM(70) <= std_logic_vector(to_signed(1013,32));
ROM(71) <= std_logic_vector(to_signed(1009,32));
ROM(72) <= std_logic_vector(to_signed(1004,32));
ROM(73) <= std_logic_vector(to_signed(999,32));
ROM(74) <= std_logic_vector(to_signed(993,32));
ROM(75) <= std_logic_vector(to_signed(987,32));
ROM(76) <= std_logic_vector(to_signed(980,32));
ROM(77) <= std_logic_vector(to_signed(972,32));
ROM(78) <= std_logic_vector(to_signed(964,32));
ROM(79) <= std_logic_vector(to_signed(955,32));
ROM(80) <= std_logic_vector(to_signed(946,32));
ROM(81) <= std_logic_vector(to_signed(936,32));
ROM(82) <= std_logic_vector(to_signed(926,32));
ROM(83) <= std_logic_vector(to_signed(915,32));
ROM(84) <= std_logic_vector(to_signed(903,32));
ROM(85) <= std_logic_vector(to_signed(891,32));
ROM(86) <= std_logic_vector(to_signed(878,32));
ROM(87) <= std_logic_vector(to_signed(865,32));
ROM(88) <= std_logic_vector(to_signed(851,32));
ROM(89) <= std_logic_vector(to_signed(837,32));
ROM(90) <= std_logic_vector(to_signed(822,32));
ROM(91) <= std_logic_vector(to_signed(807,32));
ROM(92) <= std_logic_vector(to_signed(792,32));
ROM(93) <= std_logic_vector(to_signed(775,32));
ROM(94) <= std_logic_vector(to_signed(759,32));
ROM(95) <= std_logic_vector(to_signed(742,32));
ROM(96) <= std_logic_vector(to_signed(724,32));
ROM(97) <= std_logic_vector(to_signed(706,32));
ROM(98) <= std_logic_vector(to_signed(688,32));
ROM(99) <= std_logic_vector(to_signed(669,32));
ROM(100) <= std_logic_vector(to_signed(650,32));
ROM(101) <= std_logic_vector(to_signed(630,32));
ROM(102) <= std_logic_vector(to_signed(610,32));
ROM(103) <= std_logic_vector(to_signed(590,32));
ROM(104) <= std_logic_vector(to_signed(569,32));
ROM(105) <= std_logic_vector(to_signed(548,32));
ROM(106) <= std_logic_vector(to_signed(526,32));
ROM(107) <= std_logic_vector(to_signed(505,32));
ROM(108) <= std_logic_vector(to_signed(483,32));
ROM(109) <= std_logic_vector(to_signed(460,32));
ROM(110) <= std_logic_vector(to_signed(438,32));
ROM(111) <= std_logic_vector(to_signed(415,32));
ROM(112) <= std_logic_vector(to_signed(392,32));
ROM(113) <= std_logic_vector(to_signed(369,32));
ROM(114) <= std_logic_vector(to_signed(345,32));
ROM(115) <= std_logic_vector(to_signed(321,32));
ROM(116) <= std_logic_vector(to_signed(297,32));
ROM(117) <= std_logic_vector(to_signed(273,32));
ROM(118) <= std_logic_vector(to_signed(249,32));
ROM(119) <= std_logic_vector(to_signed(224,32));
ROM(120) <= std_logic_vector(to_signed(200,32));
ROM(121) <= std_logic_vector(to_signed(175,32));
ROM(122) <= std_logic_vector(to_signed(150,32));
ROM(123) <= std_logic_vector(to_signed(125,32));
ROM(124) <= std_logic_vector(to_signed(100,32));
ROM(125) <= std_logic_vector(to_signed(75,32));
ROM(126) <= std_logic_vector(to_signed(50,32));
ROM(127) <= std_logic_vector(to_signed(25,32));
ROM(128) <= std_logic_vector(to_signed(0,32));
ROM(129) <= std_logic_vector(to_signed(-25,32));
ROM(130) <= std_logic_vector(to_signed(-50,32));
ROM(131) <= std_logic_vector(to_signed(-75,32));
ROM(132) <= std_logic_vector(to_signed(-100,32));
ROM(133) <= std_logic_vector(to_signed(-125,32));
ROM(134) <= std_logic_vector(to_signed(-150,32));
ROM(135) <= std_logic_vector(to_signed(-175,32));
ROM(136) <= std_logic_vector(to_signed(-200,32));
ROM(137) <= std_logic_vector(to_signed(-224,32));
ROM(138) <= std_logic_vector(to_signed(-249,32));
ROM(139) <= std_logic_vector(to_signed(-273,32));
ROM(140) <= std_logic_vector(to_signed(-297,32));
ROM(141) <= std_logic_vector(to_signed(-321,32));
ROM(142) <= std_logic_vector(to_signed(-345,32));
ROM(143) <= std_logic_vector(to_signed(-369,32));
ROM(144) <= std_logic_vector(to_signed(-392,32));
ROM(145) <= std_logic_vector(to_signed(-415,32));
ROM(146) <= std_logic_vector(to_signed(-438,32));
ROM(147) <= std_logic_vector(to_signed(-460,32));
ROM(148) <= std_logic_vector(to_signed(-483,32));
ROM(149) <= std_logic_vector(to_signed(-505,32));
ROM(150) <= std_logic_vector(to_signed(-526,32));
ROM(151) <= std_logic_vector(to_signed(-548,32));
ROM(152) <= std_logic_vector(to_signed(-569,32));
ROM(153) <= std_logic_vector(to_signed(-590,32));
ROM(154) <= std_logic_vector(to_signed(-610,32));
ROM(155) <= std_logic_vector(to_signed(-630,32));
ROM(156) <= std_logic_vector(to_signed(-650,32));
ROM(157) <= std_logic_vector(to_signed(-669,32));
ROM(158) <= std_logic_vector(to_signed(-688,32));
ROM(159) <= std_logic_vector(to_signed(-706,32));
ROM(160) <= std_logic_vector(to_signed(-724,32));
ROM(161) <= std_logic_vector(to_signed(-742,32));
ROM(162) <= std_logic_vector(to_signed(-759,32));
ROM(163) <= std_logic_vector(to_signed(-775,32));
ROM(164) <= std_logic_vector(to_signed(-792,32));
ROM(165) <= std_logic_vector(to_signed(-807,32));
ROM(166) <= std_logic_vector(to_signed(-822,32));
ROM(167) <= std_logic_vector(to_signed(-837,32));
ROM(168) <= std_logic_vector(to_signed(-851,32));
ROM(169) <= std_logic_vector(to_signed(-865,32));
ROM(170) <= std_logic_vector(to_signed(-878,32));
ROM(171) <= std_logic_vector(to_signed(-891,32));
ROM(172) <= std_logic_vector(to_signed(-903,32));
ROM(173) <= std_logic_vector(to_signed(-915,32));
ROM(174) <= std_logic_vector(to_signed(-926,32));
ROM(175) <= std_logic_vector(to_signed(-936,32));
ROM(176) <= std_logic_vector(to_signed(-946,32));
ROM(177) <= std_logic_vector(to_signed(-955,32));
ROM(178) <= std_logic_vector(to_signed(-964,32));
ROM(179) <= std_logic_vector(to_signed(-972,32));
ROM(180) <= std_logic_vector(to_signed(-980,32));
ROM(181) <= std_logic_vector(to_signed(-987,32));
ROM(182) <= std_logic_vector(to_signed(-993,32));
ROM(183) <= std_logic_vector(to_signed(-999,32));
ROM(184) <= std_logic_vector(to_signed(-1004,32));
ROM(185) <= std_logic_vector(to_signed(-1009,32));
ROM(186) <= std_logic_vector(to_signed(-1013,32));
ROM(187) <= std_logic_vector(to_signed(-1016,32));
ROM(188) <= std_logic_vector(to_signed(-1019,32));
ROM(189) <= std_logic_vector(to_signed(-1021,32));
ROM(190) <= std_logic_vector(to_signed(-1023,32));
ROM(191) <= std_logic_vector(to_signed(-1024,32));
ROM(192) <= std_logic_vector(to_signed(-1024,32));
ROM(193) <= std_logic_vector(to_signed(-1024,32));
ROM(194) <= std_logic_vector(to_signed(-1023,32));
ROM(195) <= std_logic_vector(to_signed(-1021,32));
ROM(196) <= std_logic_vector(to_signed(-1019,32));
ROM(197) <= std_logic_vector(to_signed(-1016,32));
ROM(198) <= std_logic_vector(to_signed(-1013,32));
ROM(199) <= std_logic_vector(to_signed(-1009,32));
ROM(200) <= std_logic_vector(to_signed(-1004,32));
ROM(201) <= std_logic_vector(to_signed(-999,32));
ROM(202) <= std_logic_vector(to_signed(-993,32));
ROM(203) <= std_logic_vector(to_signed(-987,32));
ROM(204) <= std_logic_vector(to_signed(-980,32));
ROM(205) <= std_logic_vector(to_signed(-972,32));
ROM(206) <= std_logic_vector(to_signed(-964,32));
ROM(207) <= std_logic_vector(to_signed(-955,32));
ROM(208) <= std_logic_vector(to_signed(-946,32));
ROM(209) <= std_logic_vector(to_signed(-936,32));
ROM(210) <= std_logic_vector(to_signed(-926,32));
ROM(211) <= std_logic_vector(to_signed(-915,32));
ROM(212) <= std_logic_vector(to_signed(-903,32));
ROM(213) <= std_logic_vector(to_signed(-891,32));
ROM(214) <= std_logic_vector(to_signed(-878,32));
ROM(215) <= std_logic_vector(to_signed(-865,32));
ROM(216) <= std_logic_vector(to_signed(-851,32));
ROM(217) <= std_logic_vector(to_signed(-837,32));
ROM(218) <= std_logic_vector(to_signed(-822,32));
ROM(219) <= std_logic_vector(to_signed(-807,32));
ROM(220) <= std_logic_vector(to_signed(-792,32));
ROM(221) <= std_logic_vector(to_signed(-775,32));
ROM(222) <= std_logic_vector(to_signed(-759,32));
ROM(223) <= std_logic_vector(to_signed(-742,32));
ROM(224) <= std_logic_vector(to_signed(-724,32));
ROM(225) <= std_logic_vector(to_signed(-706,32));
ROM(226) <= std_logic_vector(to_signed(-688,32));
ROM(227) <= std_logic_vector(to_signed(-669,32));
ROM(228) <= std_logic_vector(to_signed(-650,32));
ROM(229) <= std_logic_vector(to_signed(-630,32));
ROM(230) <= std_logic_vector(to_signed(-610,32));
ROM(231) <= std_logic_vector(to_signed(-590,32));
ROM(232) <= std_logic_vector(to_signed(-569,32));
ROM(233) <= std_logic_vector(to_signed(-548,32));
ROM(234) <= std_logic_vector(to_signed(-526,32));
ROM(235) <= std_logic_vector(to_signed(-505,32));
ROM(236) <= std_logic_vector(to_signed(-483,32));
ROM(237) <= std_logic_vector(to_signed(-460,32));
ROM(238) <= std_logic_vector(to_signed(-438,32));
ROM(239) <= std_logic_vector(to_signed(-415,32));
ROM(240) <= std_logic_vector(to_signed(-392,32));
ROM(241) <= std_logic_vector(to_signed(-369,32));
ROM(242) <= std_logic_vector(to_signed(-345,32));
ROM(243) <= std_logic_vector(to_signed(-321,32));
ROM(244) <= std_logic_vector(to_signed(-297,32));
ROM(245) <= std_logic_vector(to_signed(-273,32));
ROM(246) <= std_logic_vector(to_signed(-249,32));
ROM(247) <= std_logic_vector(to_signed(-224,32));
ROM(248) <= std_logic_vector(to_signed(-200,32));
ROM(249) <= std_logic_vector(to_signed(-175,32));
ROM(250) <= std_logic_vector(to_signed(-150,32));
ROM(251) <= std_logic_vector(to_signed(-125,32));
ROM(252) <= std_logic_vector(to_signed(-100,32));
ROM(253) <= std_logic_vector(to_signed(-75,32));
ROM(254) <= std_logic_vector(to_signed(-50,32));
ROM(255) <= std_logic_vector(to_signed(-25,32));
                                                                              
process(clk)                                                                  
begin                                                                         
    if rising_edge(clk) then                                                  
        if rd_en='1' then                                                   
            for I in 0 to 511 loop                                             
              if to_integer(unsigned(addr_in))=I then                         
                data_out <= ROM(I);                                           
              end if;                                                         
            end loop;                                                         
        end if;                                                               
        data_out_en <= rd_en;                                                 
    end if;                                                                   
end process;                                                                  
                                                                              
end rtl;                                                                      
