library IEEE;                                                                 
use IEEE.std_logic_1164.all;                                                  
use IEEE.numeric_std.all;                                                     
                                                                              
entity test is                                                                  
 port (                                                                       
            clk             : in std_logic;                                   
            addr_in         : in std_logic_vector(11 downto 0);               
                                                                              
            data_out        : out std_logic_vector(15 downto 0)              
 );                                                                           
end entity test;                                                                
                                                                              
architecture rtl of test is                                                     
                                                                              
type ROM_type is array (0 to 4095) of std_logic_vector(15 downto 0);            
function init_rom                                                           
	return ROM_type is                                                       
	variable tmp : ROM_type := (others => (others => '0'));                  
	begin                                                                    
        tmp(0) := std_logic_vector(to_signed(0,16));
        tmp(1) := std_logic_vector(to_signed(50,16));
        tmp(2) := std_logic_vector(to_signed(101,16));
        tmp(3) := std_logic_vector(to_signed(151,16));
        tmp(4) := std_logic_vector(to_signed(201,16));
        tmp(5) := std_logic_vector(to_signed(251,16));
        tmp(6) := std_logic_vector(to_signed(302,16));
        tmp(7) := std_logic_vector(to_signed(352,16));
        tmp(8) := std_logic_vector(to_signed(402,16));
        tmp(9) := std_logic_vector(to_signed(452,16));
        tmp(10) := std_logic_vector(to_signed(503,16));
        tmp(11) := std_logic_vector(to_signed(553,16));
        tmp(12) := std_logic_vector(to_signed(603,16));
        tmp(13) := std_logic_vector(to_signed(653,16));
        tmp(14) := std_logic_vector(to_signed(704,16));
        tmp(15) := std_logic_vector(to_signed(754,16));
        tmp(16) := std_logic_vector(to_signed(804,16));
        tmp(17) := std_logic_vector(to_signed(854,16));
        tmp(18) := std_logic_vector(to_signed(905,16));
        tmp(19) := std_logic_vector(to_signed(955,16));
        tmp(20) := std_logic_vector(to_signed(1005,16));
        tmp(21) := std_logic_vector(to_signed(1055,16));
        tmp(22) := std_logic_vector(to_signed(1106,16));
        tmp(23) := std_logic_vector(to_signed(1156,16));
        tmp(24) := std_logic_vector(to_signed(1206,16));
        tmp(25) := std_logic_vector(to_signed(1256,16));
        tmp(26) := std_logic_vector(to_signed(1307,16));
        tmp(27) := std_logic_vector(to_signed(1357,16));
        tmp(28) := std_logic_vector(to_signed(1407,16));
        tmp(29) := std_logic_vector(to_signed(1457,16));
        tmp(30) := std_logic_vector(to_signed(1507,16));
        tmp(31) := std_logic_vector(to_signed(1558,16));
        tmp(32) := std_logic_vector(to_signed(1608,16));
        tmp(33) := std_logic_vector(to_signed(1658,16));
        tmp(34) := std_logic_vector(to_signed(1708,16));
        tmp(35) := std_logic_vector(to_signed(1758,16));
        tmp(36) := std_logic_vector(to_signed(1809,16));
        tmp(37) := std_logic_vector(to_signed(1859,16));
        tmp(38) := std_logic_vector(to_signed(1909,16));
        tmp(39) := std_logic_vector(to_signed(1959,16));
        tmp(40) := std_logic_vector(to_signed(2009,16));
        tmp(41) := std_logic_vector(to_signed(2059,16));
        tmp(42) := std_logic_vector(to_signed(2110,16));
        tmp(43) := std_logic_vector(to_signed(2160,16));
        tmp(44) := std_logic_vector(to_signed(2210,16));
        tmp(45) := std_logic_vector(to_signed(2260,16));
        tmp(46) := std_logic_vector(to_signed(2310,16));
        tmp(47) := std_logic_vector(to_signed(2360,16));
        tmp(48) := std_logic_vector(to_signed(2410,16));
        tmp(49) := std_logic_vector(to_signed(2461,16));
        tmp(50) := std_logic_vector(to_signed(2511,16));
        tmp(51) := std_logic_vector(to_signed(2561,16));
        tmp(52) := std_logic_vector(to_signed(2611,16));
        tmp(53) := std_logic_vector(to_signed(2661,16));
        tmp(54) := std_logic_vector(to_signed(2711,16));
        tmp(55) := std_logic_vector(to_signed(2761,16));
        tmp(56) := std_logic_vector(to_signed(2811,16));
        tmp(57) := std_logic_vector(to_signed(2861,16));
        tmp(58) := std_logic_vector(to_signed(2911,16));
        tmp(59) := std_logic_vector(to_signed(2962,16));
        tmp(60) := std_logic_vector(to_signed(3012,16));
        tmp(61) := std_logic_vector(to_signed(3062,16));
        tmp(62) := std_logic_vector(to_signed(3112,16));
        tmp(63) := std_logic_vector(to_signed(3162,16));
        tmp(64) := std_logic_vector(to_signed(3212,16));
        tmp(65) := std_logic_vector(to_signed(3262,16));
        tmp(66) := std_logic_vector(to_signed(3312,16));
        tmp(67) := std_logic_vector(to_signed(3362,16));
        tmp(68) := std_logic_vector(to_signed(3412,16));
        tmp(69) := std_logic_vector(to_signed(3462,16));
        tmp(70) := std_logic_vector(to_signed(3512,16));
        tmp(71) := std_logic_vector(to_signed(3562,16));
        tmp(72) := std_logic_vector(to_signed(3612,16));
        tmp(73) := std_logic_vector(to_signed(3662,16));
        tmp(74) := std_logic_vector(to_signed(3712,16));
        tmp(75) := std_logic_vector(to_signed(3761,16));
        tmp(76) := std_logic_vector(to_signed(3811,16));
        tmp(77) := std_logic_vector(to_signed(3861,16));
        tmp(78) := std_logic_vector(to_signed(3911,16));
        tmp(79) := std_logic_vector(to_signed(3961,16));
        tmp(80) := std_logic_vector(to_signed(4011,16));
        tmp(81) := std_logic_vector(to_signed(4061,16));
        tmp(82) := std_logic_vector(to_signed(4111,16));
        tmp(83) := std_logic_vector(to_signed(4161,16));
        tmp(84) := std_logic_vector(to_signed(4210,16));
        tmp(85) := std_logic_vector(to_signed(4260,16));
        tmp(86) := std_logic_vector(to_signed(4310,16));
        tmp(87) := std_logic_vector(to_signed(4360,16));
        tmp(88) := std_logic_vector(to_signed(4410,16));
        tmp(89) := std_logic_vector(to_signed(4460,16));
        tmp(90) := std_logic_vector(to_signed(4509,16));
        tmp(91) := std_logic_vector(to_signed(4559,16));
        tmp(92) := std_logic_vector(to_signed(4609,16));
        tmp(93) := std_logic_vector(to_signed(4659,16));
        tmp(94) := std_logic_vector(to_signed(4708,16));
        tmp(95) := std_logic_vector(to_signed(4758,16));
        tmp(96) := std_logic_vector(to_signed(4808,16));
        tmp(97) := std_logic_vector(to_signed(4858,16));
        tmp(98) := std_logic_vector(to_signed(4907,16));
        tmp(99) := std_logic_vector(to_signed(4957,16));
        tmp(100) := std_logic_vector(to_signed(5007,16));
        tmp(101) := std_logic_vector(to_signed(5056,16));
        tmp(102) := std_logic_vector(to_signed(5106,16));
        tmp(103) := std_logic_vector(to_signed(5156,16));
        tmp(104) := std_logic_vector(to_signed(5205,16));
        tmp(105) := std_logic_vector(to_signed(5255,16));
        tmp(106) := std_logic_vector(to_signed(5305,16));
        tmp(107) := std_logic_vector(to_signed(5354,16));
        tmp(108) := std_logic_vector(to_signed(5404,16));
        tmp(109) := std_logic_vector(to_signed(5453,16));
        tmp(110) := std_logic_vector(to_signed(5503,16));
        tmp(111) := std_logic_vector(to_signed(5552,16));
        tmp(112) := std_logic_vector(to_signed(5602,16));
        tmp(113) := std_logic_vector(to_signed(5651,16));
        tmp(114) := std_logic_vector(to_signed(5701,16));
        tmp(115) := std_logic_vector(to_signed(5750,16));
        tmp(116) := std_logic_vector(to_signed(5800,16));
        tmp(117) := std_logic_vector(to_signed(5849,16));
        tmp(118) := std_logic_vector(to_signed(5899,16));
        tmp(119) := std_logic_vector(to_signed(5948,16));
        tmp(120) := std_logic_vector(to_signed(5998,16));
        tmp(121) := std_logic_vector(to_signed(6047,16));
        tmp(122) := std_logic_vector(to_signed(6096,16));
        tmp(123) := std_logic_vector(to_signed(6146,16));
        tmp(124) := std_logic_vector(to_signed(6195,16));
        tmp(125) := std_logic_vector(to_signed(6245,16));
        tmp(126) := std_logic_vector(to_signed(6294,16));
        tmp(127) := std_logic_vector(to_signed(6343,16));
        tmp(128) := std_logic_vector(to_signed(6393,16));
        tmp(129) := std_logic_vector(to_signed(6442,16));
        tmp(130) := std_logic_vector(to_signed(6491,16));
        tmp(131) := std_logic_vector(to_signed(6540,16));
        tmp(132) := std_logic_vector(to_signed(6590,16));
        tmp(133) := std_logic_vector(to_signed(6639,16));
        tmp(134) := std_logic_vector(to_signed(6688,16));
        tmp(135) := std_logic_vector(to_signed(6737,16));
        tmp(136) := std_logic_vector(to_signed(6786,16));
        tmp(137) := std_logic_vector(to_signed(6836,16));
        tmp(138) := std_logic_vector(to_signed(6885,16));
        tmp(139) := std_logic_vector(to_signed(6934,16));
        tmp(140) := std_logic_vector(to_signed(6983,16));
        tmp(141) := std_logic_vector(to_signed(7032,16));
        tmp(142) := std_logic_vector(to_signed(7081,16));
        tmp(143) := std_logic_vector(to_signed(7130,16));
        tmp(144) := std_logic_vector(to_signed(7179,16));
        tmp(145) := std_logic_vector(to_signed(7228,16));
        tmp(146) := std_logic_vector(to_signed(7277,16));
        tmp(147) := std_logic_vector(to_signed(7326,16));
        tmp(148) := std_logic_vector(to_signed(7375,16));
        tmp(149) := std_logic_vector(to_signed(7424,16));
        tmp(150) := std_logic_vector(to_signed(7473,16));
        tmp(151) := std_logic_vector(to_signed(7522,16));
        tmp(152) := std_logic_vector(to_signed(7571,16));
        tmp(153) := std_logic_vector(to_signed(7620,16));
        tmp(154) := std_logic_vector(to_signed(7669,16));
        tmp(155) := std_logic_vector(to_signed(7718,16));
        tmp(156) := std_logic_vector(to_signed(7767,16));
        tmp(157) := std_logic_vector(to_signed(7815,16));
        tmp(158) := std_logic_vector(to_signed(7864,16));
        tmp(159) := std_logic_vector(to_signed(7913,16));
        tmp(160) := std_logic_vector(to_signed(7962,16));
        tmp(161) := std_logic_vector(to_signed(8010,16));
        tmp(162) := std_logic_vector(to_signed(8059,16));
        tmp(163) := std_logic_vector(to_signed(8108,16));
        tmp(164) := std_logic_vector(to_signed(8157,16));
        tmp(165) := std_logic_vector(to_signed(8205,16));
        tmp(166) := std_logic_vector(to_signed(8254,16));
        tmp(167) := std_logic_vector(to_signed(8303,16));
        tmp(168) := std_logic_vector(to_signed(8351,16));
        tmp(169) := std_logic_vector(to_signed(8400,16));
        tmp(170) := std_logic_vector(to_signed(8448,16));
        tmp(171) := std_logic_vector(to_signed(8497,16));
        tmp(172) := std_logic_vector(to_signed(8545,16));
        tmp(173) := std_logic_vector(to_signed(8594,16));
        tmp(174) := std_logic_vector(to_signed(8642,16));
        tmp(175) := std_logic_vector(to_signed(8691,16));
        tmp(176) := std_logic_vector(to_signed(8739,16));
        tmp(177) := std_logic_vector(to_signed(8788,16));
        tmp(178) := std_logic_vector(to_signed(8836,16));
        tmp(179) := std_logic_vector(to_signed(8885,16));
        tmp(180) := std_logic_vector(to_signed(8933,16));
        tmp(181) := std_logic_vector(to_signed(8981,16));
        tmp(182) := std_logic_vector(to_signed(9030,16));
        tmp(183) := std_logic_vector(to_signed(9078,16));
        tmp(184) := std_logic_vector(to_signed(9126,16));
        tmp(185) := std_logic_vector(to_signed(9175,16));
        tmp(186) := std_logic_vector(to_signed(9223,16));
        tmp(187) := std_logic_vector(to_signed(9271,16));
        tmp(188) := std_logic_vector(to_signed(9319,16));
        tmp(189) := std_logic_vector(to_signed(9367,16));
        tmp(190) := std_logic_vector(to_signed(9416,16));
        tmp(191) := std_logic_vector(to_signed(9464,16));
        tmp(192) := std_logic_vector(to_signed(9512,16));
        tmp(193) := std_logic_vector(to_signed(9560,16));
        tmp(194) := std_logic_vector(to_signed(9608,16));
        tmp(195) := std_logic_vector(to_signed(9656,16));
        tmp(196) := std_logic_vector(to_signed(9704,16));
        tmp(197) := std_logic_vector(to_signed(9752,16));
        tmp(198) := std_logic_vector(to_signed(9800,16));
        tmp(199) := std_logic_vector(to_signed(9848,16));
        tmp(200) := std_logic_vector(to_signed(9896,16));
        tmp(201) := std_logic_vector(to_signed(9944,16));
        tmp(202) := std_logic_vector(to_signed(9992,16));
        tmp(203) := std_logic_vector(to_signed(10039,16));
        tmp(204) := std_logic_vector(to_signed(10087,16));
        tmp(205) := std_logic_vector(to_signed(10135,16));
        tmp(206) := std_logic_vector(to_signed(10183,16));
        tmp(207) := std_logic_vector(to_signed(10231,16));
        tmp(208) := std_logic_vector(to_signed(10278,16));
        tmp(209) := std_logic_vector(to_signed(10326,16));
        tmp(210) := std_logic_vector(to_signed(10374,16));
        tmp(211) := std_logic_vector(to_signed(10421,16));
        tmp(212) := std_logic_vector(to_signed(10469,16));
        tmp(213) := std_logic_vector(to_signed(10517,16));
        tmp(214) := std_logic_vector(to_signed(10564,16));
        tmp(215) := std_logic_vector(to_signed(10612,16));
        tmp(216) := std_logic_vector(to_signed(10659,16));
        tmp(217) := std_logic_vector(to_signed(10707,16));
        tmp(218) := std_logic_vector(to_signed(10754,16));
        tmp(219) := std_logic_vector(to_signed(10802,16));
        tmp(220) := std_logic_vector(to_signed(10849,16));
        tmp(221) := std_logic_vector(to_signed(10897,16));
        tmp(222) := std_logic_vector(to_signed(10944,16));
        tmp(223) := std_logic_vector(to_signed(10992,16));
        tmp(224) := std_logic_vector(to_signed(11039,16));
        tmp(225) := std_logic_vector(to_signed(11086,16));
        tmp(226) := std_logic_vector(to_signed(11133,16));
        tmp(227) := std_logic_vector(to_signed(11181,16));
        tmp(228) := std_logic_vector(to_signed(11228,16));
        tmp(229) := std_logic_vector(to_signed(11275,16));
        tmp(230) := std_logic_vector(to_signed(11322,16));
        tmp(231) := std_logic_vector(to_signed(11370,16));
        tmp(232) := std_logic_vector(to_signed(11417,16));
        tmp(233) := std_logic_vector(to_signed(11464,16));
        tmp(234) := std_logic_vector(to_signed(11511,16));
        tmp(235) := std_logic_vector(to_signed(11558,16));
        tmp(236) := std_logic_vector(to_signed(11605,16));
        tmp(237) := std_logic_vector(to_signed(11652,16));
        tmp(238) := std_logic_vector(to_signed(11699,16));
        tmp(239) := std_logic_vector(to_signed(11746,16));
        tmp(240) := std_logic_vector(to_signed(11793,16));
        tmp(241) := std_logic_vector(to_signed(11840,16));
        tmp(242) := std_logic_vector(to_signed(11886,16));
        tmp(243) := std_logic_vector(to_signed(11933,16));
        tmp(244) := std_logic_vector(to_signed(11980,16));
        tmp(245) := std_logic_vector(to_signed(12027,16));
        tmp(246) := std_logic_vector(to_signed(12074,16));
        tmp(247) := std_logic_vector(to_signed(12120,16));
        tmp(248) := std_logic_vector(to_signed(12167,16));
        tmp(249) := std_logic_vector(to_signed(12214,16));
        tmp(250) := std_logic_vector(to_signed(12260,16));
        tmp(251) := std_logic_vector(to_signed(12307,16));
        tmp(252) := std_logic_vector(to_signed(12353,16));
        tmp(253) := std_logic_vector(to_signed(12400,16));
        tmp(254) := std_logic_vector(to_signed(12446,16));
        tmp(255) := std_logic_vector(to_signed(12493,16));
        tmp(256) := std_logic_vector(to_signed(12539,16));
        tmp(257) := std_logic_vector(to_signed(12586,16));
        tmp(258) := std_logic_vector(to_signed(12632,16));
        tmp(259) := std_logic_vector(to_signed(12679,16));
        tmp(260) := std_logic_vector(to_signed(12725,16));
        tmp(261) := std_logic_vector(to_signed(12771,16));
        tmp(262) := std_logic_vector(to_signed(12817,16));
        tmp(263) := std_logic_vector(to_signed(12864,16));
        tmp(264) := std_logic_vector(to_signed(12910,16));
        tmp(265) := std_logic_vector(to_signed(12956,16));
        tmp(266) := std_logic_vector(to_signed(13002,16));
        tmp(267) := std_logic_vector(to_signed(13048,16));
        tmp(268) := std_logic_vector(to_signed(13094,16));
        tmp(269) := std_logic_vector(to_signed(13141,16));
        tmp(270) := std_logic_vector(to_signed(13187,16));
        tmp(271) := std_logic_vector(to_signed(13233,16));
        tmp(272) := std_logic_vector(to_signed(13279,16));
        tmp(273) := std_logic_vector(to_signed(13324,16));
        tmp(274) := std_logic_vector(to_signed(13370,16));
        tmp(275) := std_logic_vector(to_signed(13416,16));
        tmp(276) := std_logic_vector(to_signed(13462,16));
        tmp(277) := std_logic_vector(to_signed(13508,16));
        tmp(278) := std_logic_vector(to_signed(13554,16));
        tmp(279) := std_logic_vector(to_signed(13599,16));
        tmp(280) := std_logic_vector(to_signed(13645,16));
        tmp(281) := std_logic_vector(to_signed(13691,16));
        tmp(282) := std_logic_vector(to_signed(13736,16));
        tmp(283) := std_logic_vector(to_signed(13782,16));
        tmp(284) := std_logic_vector(to_signed(13828,16));
        tmp(285) := std_logic_vector(to_signed(13873,16));
        tmp(286) := std_logic_vector(to_signed(13919,16));
        tmp(287) := std_logic_vector(to_signed(13964,16));
        tmp(288) := std_logic_vector(to_signed(14010,16));
        tmp(289) := std_logic_vector(to_signed(14055,16));
        tmp(290) := std_logic_vector(to_signed(14101,16));
        tmp(291) := std_logic_vector(to_signed(14146,16));
        tmp(292) := std_logic_vector(to_signed(14191,16));
        tmp(293) := std_logic_vector(to_signed(14236,16));
        tmp(294) := std_logic_vector(to_signed(14282,16));
        tmp(295) := std_logic_vector(to_signed(14327,16));
        tmp(296) := std_logic_vector(to_signed(14372,16));
        tmp(297) := std_logic_vector(to_signed(14417,16));
        tmp(298) := std_logic_vector(to_signed(14462,16));
        tmp(299) := std_logic_vector(to_signed(14507,16));
        tmp(300) := std_logic_vector(to_signed(14553,16));
        tmp(301) := std_logic_vector(to_signed(14598,16));
        tmp(302) := std_logic_vector(to_signed(14643,16));
        tmp(303) := std_logic_vector(to_signed(14688,16));
        tmp(304) := std_logic_vector(to_signed(14732,16));
        tmp(305) := std_logic_vector(to_signed(14777,16));
        tmp(306) := std_logic_vector(to_signed(14822,16));
        tmp(307) := std_logic_vector(to_signed(14867,16));
        tmp(308) := std_logic_vector(to_signed(14912,16));
        tmp(309) := std_logic_vector(to_signed(14956,16));
        tmp(310) := std_logic_vector(to_signed(15001,16));
        tmp(311) := std_logic_vector(to_signed(15046,16));
        tmp(312) := std_logic_vector(to_signed(15090,16));
        tmp(313) := std_logic_vector(to_signed(15135,16));
        tmp(314) := std_logic_vector(to_signed(15180,16));
        tmp(315) := std_logic_vector(to_signed(15224,16));
        tmp(316) := std_logic_vector(to_signed(15269,16));
        tmp(317) := std_logic_vector(to_signed(15313,16));
        tmp(318) := std_logic_vector(to_signed(15358,16));
        tmp(319) := std_logic_vector(to_signed(15402,16));
        tmp(320) := std_logic_vector(to_signed(15446,16));
        tmp(321) := std_logic_vector(to_signed(15491,16));
        tmp(322) := std_logic_vector(to_signed(15535,16));
        tmp(323) := std_logic_vector(to_signed(15579,16));
        tmp(324) := std_logic_vector(to_signed(15623,16));
        tmp(325) := std_logic_vector(to_signed(15667,16));
        tmp(326) := std_logic_vector(to_signed(15712,16));
        tmp(327) := std_logic_vector(to_signed(15756,16));
        tmp(328) := std_logic_vector(to_signed(15800,16));
        tmp(329) := std_logic_vector(to_signed(15844,16));
        tmp(330) := std_logic_vector(to_signed(15888,16));
        tmp(331) := std_logic_vector(to_signed(15932,16));
        tmp(332) := std_logic_vector(to_signed(15976,16));
        tmp(333) := std_logic_vector(to_signed(16019,16));
        tmp(334) := std_logic_vector(to_signed(16063,16));
        tmp(335) := std_logic_vector(to_signed(16107,16));
        tmp(336) := std_logic_vector(to_signed(16151,16));
        tmp(337) := std_logic_vector(to_signed(16195,16));
        tmp(338) := std_logic_vector(to_signed(16238,16));
        tmp(339) := std_logic_vector(to_signed(16282,16));
        tmp(340) := std_logic_vector(to_signed(16325,16));
        tmp(341) := std_logic_vector(to_signed(16369,16));
        tmp(342) := std_logic_vector(to_signed(16413,16));
        tmp(343) := std_logic_vector(to_signed(16456,16));
        tmp(344) := std_logic_vector(to_signed(16499,16));
        tmp(345) := std_logic_vector(to_signed(16543,16));
        tmp(346) := std_logic_vector(to_signed(16586,16));
        tmp(347) := std_logic_vector(to_signed(16630,16));
        tmp(348) := std_logic_vector(to_signed(16673,16));
        tmp(349) := std_logic_vector(to_signed(16716,16));
        tmp(350) := std_logic_vector(to_signed(16759,16));
        tmp(351) := std_logic_vector(to_signed(16802,16));
        tmp(352) := std_logic_vector(to_signed(16846,16));
        tmp(353) := std_logic_vector(to_signed(16889,16));
        tmp(354) := std_logic_vector(to_signed(16932,16));
        tmp(355) := std_logic_vector(to_signed(16975,16));
        tmp(356) := std_logic_vector(to_signed(17018,16));
        tmp(357) := std_logic_vector(to_signed(17061,16));
        tmp(358) := std_logic_vector(to_signed(17104,16));
        tmp(359) := std_logic_vector(to_signed(17146,16));
        tmp(360) := std_logic_vector(to_signed(17189,16));
        tmp(361) := std_logic_vector(to_signed(17232,16));
        tmp(362) := std_logic_vector(to_signed(17275,16));
        tmp(363) := std_logic_vector(to_signed(17317,16));
        tmp(364) := std_logic_vector(to_signed(17360,16));
        tmp(365) := std_logic_vector(to_signed(17403,16));
        tmp(366) := std_logic_vector(to_signed(17445,16));
        tmp(367) := std_logic_vector(to_signed(17488,16));
        tmp(368) := std_logic_vector(to_signed(17530,16));
        tmp(369) := std_logic_vector(to_signed(17573,16));
        tmp(370) := std_logic_vector(to_signed(17615,16));
        tmp(371) := std_logic_vector(to_signed(17657,16));
        tmp(372) := std_logic_vector(to_signed(17700,16));
        tmp(373) := std_logic_vector(to_signed(17742,16));
        tmp(374) := std_logic_vector(to_signed(17784,16));
        tmp(375) := std_logic_vector(to_signed(17827,16));
        tmp(376) := std_logic_vector(to_signed(17869,16));
        tmp(377) := std_logic_vector(to_signed(17911,16));
        tmp(378) := std_logic_vector(to_signed(17953,16));
        tmp(379) := std_logic_vector(to_signed(17995,16));
        tmp(380) := std_logic_vector(to_signed(18037,16));
        tmp(381) := std_logic_vector(to_signed(18079,16));
        tmp(382) := std_logic_vector(to_signed(18121,16));
        tmp(383) := std_logic_vector(to_signed(18163,16));
        tmp(384) := std_logic_vector(to_signed(18204,16));
        tmp(385) := std_logic_vector(to_signed(18246,16));
        tmp(386) := std_logic_vector(to_signed(18288,16));
        tmp(387) := std_logic_vector(to_signed(18330,16));
        tmp(388) := std_logic_vector(to_signed(18371,16));
        tmp(389) := std_logic_vector(to_signed(18413,16));
        tmp(390) := std_logic_vector(to_signed(18454,16));
        tmp(391) := std_logic_vector(to_signed(18496,16));
        tmp(392) := std_logic_vector(to_signed(18537,16));
        tmp(393) := std_logic_vector(to_signed(18579,16));
        tmp(394) := std_logic_vector(to_signed(18620,16));
        tmp(395) := std_logic_vector(to_signed(18661,16));
        tmp(396) := std_logic_vector(to_signed(18703,16));
        tmp(397) := std_logic_vector(to_signed(18744,16));
        tmp(398) := std_logic_vector(to_signed(18785,16));
        tmp(399) := std_logic_vector(to_signed(18826,16));
        tmp(400) := std_logic_vector(to_signed(18868,16));
        tmp(401) := std_logic_vector(to_signed(18909,16));
        tmp(402) := std_logic_vector(to_signed(18950,16));
        tmp(403) := std_logic_vector(to_signed(18991,16));
        tmp(404) := std_logic_vector(to_signed(19032,16));
        tmp(405) := std_logic_vector(to_signed(19072,16));
        tmp(406) := std_logic_vector(to_signed(19113,16));
        tmp(407) := std_logic_vector(to_signed(19154,16));
        tmp(408) := std_logic_vector(to_signed(19195,16));
        tmp(409) := std_logic_vector(to_signed(19236,16));
        tmp(410) := std_logic_vector(to_signed(19276,16));
        tmp(411) := std_logic_vector(to_signed(19317,16));
        tmp(412) := std_logic_vector(to_signed(19357,16));
        tmp(413) := std_logic_vector(to_signed(19398,16));
        tmp(414) := std_logic_vector(to_signed(19438,16));
        tmp(415) := std_logic_vector(to_signed(19479,16));
        tmp(416) := std_logic_vector(to_signed(19519,16));
        tmp(417) := std_logic_vector(to_signed(19560,16));
        tmp(418) := std_logic_vector(to_signed(19600,16));
        tmp(419) := std_logic_vector(to_signed(19640,16));
        tmp(420) := std_logic_vector(to_signed(19680,16));
        tmp(421) := std_logic_vector(to_signed(19721,16));
        tmp(422) := std_logic_vector(to_signed(19761,16));
        tmp(423) := std_logic_vector(to_signed(19801,16));
        tmp(424) := std_logic_vector(to_signed(19841,16));
        tmp(425) := std_logic_vector(to_signed(19881,16));
        tmp(426) := std_logic_vector(to_signed(19921,16));
        tmp(427) := std_logic_vector(to_signed(19961,16));
        tmp(428) := std_logic_vector(to_signed(20000,16));
        tmp(429) := std_logic_vector(to_signed(20040,16));
        tmp(430) := std_logic_vector(to_signed(20080,16));
        tmp(431) := std_logic_vector(to_signed(20120,16));
        tmp(432) := std_logic_vector(to_signed(20159,16));
        tmp(433) := std_logic_vector(to_signed(20199,16));
        tmp(434) := std_logic_vector(to_signed(20238,16));
        tmp(435) := std_logic_vector(to_signed(20278,16));
        tmp(436) := std_logic_vector(to_signed(20317,16));
        tmp(437) := std_logic_vector(to_signed(20357,16));
        tmp(438) := std_logic_vector(to_signed(20396,16));
        tmp(439) := std_logic_vector(to_signed(20436,16));
        tmp(440) := std_logic_vector(to_signed(20475,16));
        tmp(441) := std_logic_vector(to_signed(20514,16));
        tmp(442) := std_logic_vector(to_signed(20553,16));
        tmp(443) := std_logic_vector(to_signed(20592,16));
        tmp(444) := std_logic_vector(to_signed(20631,16));
        tmp(445) := std_logic_vector(to_signed(20670,16));
        tmp(446) := std_logic_vector(to_signed(20709,16));
        tmp(447) := std_logic_vector(to_signed(20748,16));
        tmp(448) := std_logic_vector(to_signed(20787,16));
        tmp(449) := std_logic_vector(to_signed(20826,16));
        tmp(450) := std_logic_vector(to_signed(20865,16));
        tmp(451) := std_logic_vector(to_signed(20904,16));
        tmp(452) := std_logic_vector(to_signed(20942,16));
        tmp(453) := std_logic_vector(to_signed(20981,16));
        tmp(454) := std_logic_vector(to_signed(21019,16));
        tmp(455) := std_logic_vector(to_signed(21058,16));
        tmp(456) := std_logic_vector(to_signed(21096,16));
        tmp(457) := std_logic_vector(to_signed(21135,16));
        tmp(458) := std_logic_vector(to_signed(21173,16));
        tmp(459) := std_logic_vector(to_signed(21212,16));
        tmp(460) := std_logic_vector(to_signed(21250,16));
        tmp(461) := std_logic_vector(to_signed(21288,16));
        tmp(462) := std_logic_vector(to_signed(21326,16));
        tmp(463) := std_logic_vector(to_signed(21364,16));
        tmp(464) := std_logic_vector(to_signed(21403,16));
        tmp(465) := std_logic_vector(to_signed(21441,16));
        tmp(466) := std_logic_vector(to_signed(21479,16));
        tmp(467) := std_logic_vector(to_signed(21516,16));
        tmp(468) := std_logic_vector(to_signed(21554,16));
        tmp(469) := std_logic_vector(to_signed(21592,16));
        tmp(470) := std_logic_vector(to_signed(21630,16));
        tmp(471) := std_logic_vector(to_signed(21668,16));
        tmp(472) := std_logic_vector(to_signed(21705,16));
        tmp(473) := std_logic_vector(to_signed(21743,16));
        tmp(474) := std_logic_vector(to_signed(21781,16));
        tmp(475) := std_logic_vector(to_signed(21818,16));
        tmp(476) := std_logic_vector(to_signed(21856,16));
        tmp(477) := std_logic_vector(to_signed(21893,16));
        tmp(478) := std_logic_vector(to_signed(21930,16));
        tmp(479) := std_logic_vector(to_signed(21968,16));
        tmp(480) := std_logic_vector(to_signed(22005,16));
        tmp(481) := std_logic_vector(to_signed(22042,16));
        tmp(482) := std_logic_vector(to_signed(22079,16));
        tmp(483) := std_logic_vector(to_signed(22116,16));
        tmp(484) := std_logic_vector(to_signed(22154,16));
        tmp(485) := std_logic_vector(to_signed(22191,16));
        tmp(486) := std_logic_vector(to_signed(22227,16));
        tmp(487) := std_logic_vector(to_signed(22264,16));
        tmp(488) := std_logic_vector(to_signed(22301,16));
        tmp(489) := std_logic_vector(to_signed(22338,16));
        tmp(490) := std_logic_vector(to_signed(22375,16));
        tmp(491) := std_logic_vector(to_signed(22411,16));
        tmp(492) := std_logic_vector(to_signed(22448,16));
        tmp(493) := std_logic_vector(to_signed(22485,16));
        tmp(494) := std_logic_vector(to_signed(22521,16));
        tmp(495) := std_logic_vector(to_signed(22558,16));
        tmp(496) := std_logic_vector(to_signed(22594,16));
        tmp(497) := std_logic_vector(to_signed(22631,16));
        tmp(498) := std_logic_vector(to_signed(22667,16));
        tmp(499) := std_logic_vector(to_signed(22703,16));
        tmp(500) := std_logic_vector(to_signed(22739,16));
        tmp(501) := std_logic_vector(to_signed(22776,16));
        tmp(502) := std_logic_vector(to_signed(22812,16));
        tmp(503) := std_logic_vector(to_signed(22848,16));
        tmp(504) := std_logic_vector(to_signed(22884,16));
        tmp(505) := std_logic_vector(to_signed(22920,16));
        tmp(506) := std_logic_vector(to_signed(22956,16));
        tmp(507) := std_logic_vector(to_signed(22991,16));
        tmp(508) := std_logic_vector(to_signed(23027,16));
        tmp(509) := std_logic_vector(to_signed(23063,16));
        tmp(510) := std_logic_vector(to_signed(23099,16));
        tmp(511) := std_logic_vector(to_signed(23134,16));
        tmp(512) := std_logic_vector(to_signed(23170,16));
        tmp(513) := std_logic_vector(to_signed(23205,16));
        tmp(514) := std_logic_vector(to_signed(23241,16));
        tmp(515) := std_logic_vector(to_signed(23276,16));
        tmp(516) := std_logic_vector(to_signed(23311,16));
        tmp(517) := std_logic_vector(to_signed(23347,16));
        tmp(518) := std_logic_vector(to_signed(23382,16));
        tmp(519) := std_logic_vector(to_signed(23417,16));
        tmp(520) := std_logic_vector(to_signed(23452,16));
        tmp(521) := std_logic_vector(to_signed(23487,16));
        tmp(522) := std_logic_vector(to_signed(23522,16));
        tmp(523) := std_logic_vector(to_signed(23557,16));
        tmp(524) := std_logic_vector(to_signed(23592,16));
        tmp(525) := std_logic_vector(to_signed(23627,16));
        tmp(526) := std_logic_vector(to_signed(23662,16));
        tmp(527) := std_logic_vector(to_signed(23697,16));
        tmp(528) := std_logic_vector(to_signed(23731,16));
        tmp(529) := std_logic_vector(to_signed(23766,16));
        tmp(530) := std_logic_vector(to_signed(23801,16));
        tmp(531) := std_logic_vector(to_signed(23835,16));
        tmp(532) := std_logic_vector(to_signed(23870,16));
        tmp(533) := std_logic_vector(to_signed(23904,16));
        tmp(534) := std_logic_vector(to_signed(23938,16));
        tmp(535) := std_logic_vector(to_signed(23973,16));
        tmp(536) := std_logic_vector(to_signed(24007,16));
        tmp(537) := std_logic_vector(to_signed(24041,16));
        tmp(538) := std_logic_vector(to_signed(24075,16));
        tmp(539) := std_logic_vector(to_signed(24109,16));
        tmp(540) := std_logic_vector(to_signed(24143,16));
        tmp(541) := std_logic_vector(to_signed(24177,16));
        tmp(542) := std_logic_vector(to_signed(24211,16));
        tmp(543) := std_logic_vector(to_signed(24245,16));
        tmp(544) := std_logic_vector(to_signed(24279,16));
        tmp(545) := std_logic_vector(to_signed(24312,16));
        tmp(546) := std_logic_vector(to_signed(24346,16));
        tmp(547) := std_logic_vector(to_signed(24380,16));
        tmp(548) := std_logic_vector(to_signed(24413,16));
        tmp(549) := std_logic_vector(to_signed(24447,16));
        tmp(550) := std_logic_vector(to_signed(24480,16));
        tmp(551) := std_logic_vector(to_signed(24514,16));
        tmp(552) := std_logic_vector(to_signed(24547,16));
        tmp(553) := std_logic_vector(to_signed(24580,16));
        tmp(554) := std_logic_vector(to_signed(24613,16));
        tmp(555) := std_logic_vector(to_signed(24647,16));
        tmp(556) := std_logic_vector(to_signed(24680,16));
        tmp(557) := std_logic_vector(to_signed(24713,16));
        tmp(558) := std_logic_vector(to_signed(24746,16));
        tmp(559) := std_logic_vector(to_signed(24779,16));
        tmp(560) := std_logic_vector(to_signed(24811,16));
        tmp(561) := std_logic_vector(to_signed(24844,16));
        tmp(562) := std_logic_vector(to_signed(24877,16));
        tmp(563) := std_logic_vector(to_signed(24910,16));
        tmp(564) := std_logic_vector(to_signed(24942,16));
        tmp(565) := std_logic_vector(to_signed(24975,16));
        tmp(566) := std_logic_vector(to_signed(25007,16));
        tmp(567) := std_logic_vector(to_signed(25040,16));
        tmp(568) := std_logic_vector(to_signed(25072,16));
        tmp(569) := std_logic_vector(to_signed(25105,16));
        tmp(570) := std_logic_vector(to_signed(25137,16));
        tmp(571) := std_logic_vector(to_signed(25169,16));
        tmp(572) := std_logic_vector(to_signed(25201,16));
        tmp(573) := std_logic_vector(to_signed(25233,16));
        tmp(574) := std_logic_vector(to_signed(25265,16));
        tmp(575) := std_logic_vector(to_signed(25297,16));
        tmp(576) := std_logic_vector(to_signed(25329,16));
        tmp(577) := std_logic_vector(to_signed(25361,16));
        tmp(578) := std_logic_vector(to_signed(25393,16));
        tmp(579) := std_logic_vector(to_signed(25425,16));
        tmp(580) := std_logic_vector(to_signed(25456,16));
        tmp(581) := std_logic_vector(to_signed(25488,16));
        tmp(582) := std_logic_vector(to_signed(25519,16));
        tmp(583) := std_logic_vector(to_signed(25551,16));
        tmp(584) := std_logic_vector(to_signed(25582,16));
        tmp(585) := std_logic_vector(to_signed(25614,16));
        tmp(586) := std_logic_vector(to_signed(25645,16));
        tmp(587) := std_logic_vector(to_signed(25676,16));
        tmp(588) := std_logic_vector(to_signed(25708,16));
        tmp(589) := std_logic_vector(to_signed(25739,16));
        tmp(590) := std_logic_vector(to_signed(25770,16));
        tmp(591) := std_logic_vector(to_signed(25801,16));
        tmp(592) := std_logic_vector(to_signed(25832,16));
        tmp(593) := std_logic_vector(to_signed(25863,16));
        tmp(594) := std_logic_vector(to_signed(25893,16));
        tmp(595) := std_logic_vector(to_signed(25924,16));
        tmp(596) := std_logic_vector(to_signed(25955,16));
        tmp(597) := std_logic_vector(to_signed(25986,16));
        tmp(598) := std_logic_vector(to_signed(26016,16));
        tmp(599) := std_logic_vector(to_signed(26047,16));
        tmp(600) := std_logic_vector(to_signed(26077,16));
        tmp(601) := std_logic_vector(to_signed(26108,16));
        tmp(602) := std_logic_vector(to_signed(26138,16));
        tmp(603) := std_logic_vector(to_signed(26168,16));
        tmp(604) := std_logic_vector(to_signed(26198,16));
        tmp(605) := std_logic_vector(to_signed(26229,16));
        tmp(606) := std_logic_vector(to_signed(26259,16));
        tmp(607) := std_logic_vector(to_signed(26289,16));
        tmp(608) := std_logic_vector(to_signed(26319,16));
        tmp(609) := std_logic_vector(to_signed(26349,16));
        tmp(610) := std_logic_vector(to_signed(26378,16));
        tmp(611) := std_logic_vector(to_signed(26408,16));
        tmp(612) := std_logic_vector(to_signed(26438,16));
        tmp(613) := std_logic_vector(to_signed(26468,16));
        tmp(614) := std_logic_vector(to_signed(26497,16));
        tmp(615) := std_logic_vector(to_signed(26527,16));
        tmp(616) := std_logic_vector(to_signed(26556,16));
        tmp(617) := std_logic_vector(to_signed(26586,16));
        tmp(618) := std_logic_vector(to_signed(26615,16));
        tmp(619) := std_logic_vector(to_signed(26644,16));
        tmp(620) := std_logic_vector(to_signed(26674,16));
        tmp(621) := std_logic_vector(to_signed(26703,16));
        tmp(622) := std_logic_vector(to_signed(26732,16));
        tmp(623) := std_logic_vector(to_signed(26761,16));
        tmp(624) := std_logic_vector(to_signed(26790,16));
        tmp(625) := std_logic_vector(to_signed(26819,16));
        tmp(626) := std_logic_vector(to_signed(26848,16));
        tmp(627) := std_logic_vector(to_signed(26876,16));
        tmp(628) := std_logic_vector(to_signed(26905,16));
        tmp(629) := std_logic_vector(to_signed(26934,16));
        tmp(630) := std_logic_vector(to_signed(26962,16));
        tmp(631) := std_logic_vector(to_signed(26991,16));
        tmp(632) := std_logic_vector(to_signed(27019,16));
        tmp(633) := std_logic_vector(to_signed(27048,16));
        tmp(634) := std_logic_vector(to_signed(27076,16));
        tmp(635) := std_logic_vector(to_signed(27104,16));
        tmp(636) := std_logic_vector(to_signed(27133,16));
        tmp(637) := std_logic_vector(to_signed(27161,16));
        tmp(638) := std_logic_vector(to_signed(27189,16));
        tmp(639) := std_logic_vector(to_signed(27217,16));
        tmp(640) := std_logic_vector(to_signed(27245,16));
        tmp(641) := std_logic_vector(to_signed(27273,16));
        tmp(642) := std_logic_vector(to_signed(27300,16));
        tmp(643) := std_logic_vector(to_signed(27328,16));
        tmp(644) := std_logic_vector(to_signed(27356,16));
        tmp(645) := std_logic_vector(to_signed(27384,16));
        tmp(646) := std_logic_vector(to_signed(27411,16));
        tmp(647) := std_logic_vector(to_signed(27439,16));
        tmp(648) := std_logic_vector(to_signed(27466,16));
        tmp(649) := std_logic_vector(to_signed(27493,16));
        tmp(650) := std_logic_vector(to_signed(27521,16));
        tmp(651) := std_logic_vector(to_signed(27548,16));
        tmp(652) := std_logic_vector(to_signed(27575,16));
        tmp(653) := std_logic_vector(to_signed(27602,16));
        tmp(654) := std_logic_vector(to_signed(27629,16));
        tmp(655) := std_logic_vector(to_signed(27656,16));
        tmp(656) := std_logic_vector(to_signed(27683,16));
        tmp(657) := std_logic_vector(to_signed(27710,16));
        tmp(658) := std_logic_vector(to_signed(27737,16));
        tmp(659) := std_logic_vector(to_signed(27764,16));
        tmp(660) := std_logic_vector(to_signed(27790,16));
        tmp(661) := std_logic_vector(to_signed(27817,16));
        tmp(662) := std_logic_vector(to_signed(27843,16));
        tmp(663) := std_logic_vector(to_signed(27870,16));
        tmp(664) := std_logic_vector(to_signed(27896,16));
        tmp(665) := std_logic_vector(to_signed(27923,16));
        tmp(666) := std_logic_vector(to_signed(27949,16));
        tmp(667) := std_logic_vector(to_signed(27975,16));
        tmp(668) := std_logic_vector(to_signed(28001,16));
        tmp(669) := std_logic_vector(to_signed(28027,16));
        tmp(670) := std_logic_vector(to_signed(28053,16));
        tmp(671) := std_logic_vector(to_signed(28079,16));
        tmp(672) := std_logic_vector(to_signed(28105,16));
        tmp(673) := std_logic_vector(to_signed(28131,16));
        tmp(674) := std_logic_vector(to_signed(28157,16));
        tmp(675) := std_logic_vector(to_signed(28182,16));
        tmp(676) := std_logic_vector(to_signed(28208,16));
        tmp(677) := std_logic_vector(to_signed(28234,16));
        tmp(678) := std_logic_vector(to_signed(28259,16));
        tmp(679) := std_logic_vector(to_signed(28284,16));
        tmp(680) := std_logic_vector(to_signed(28310,16));
        tmp(681) := std_logic_vector(to_signed(28335,16));
        tmp(682) := std_logic_vector(to_signed(28360,16));
        tmp(683) := std_logic_vector(to_signed(28385,16));
        tmp(684) := std_logic_vector(to_signed(28411,16));
        tmp(685) := std_logic_vector(to_signed(28436,16));
        tmp(686) := std_logic_vector(to_signed(28460,16));
        tmp(687) := std_logic_vector(to_signed(28485,16));
        tmp(688) := std_logic_vector(to_signed(28510,16));
        tmp(689) := std_logic_vector(to_signed(28535,16));
        tmp(690) := std_logic_vector(to_signed(28560,16));
        tmp(691) := std_logic_vector(to_signed(28584,16));
        tmp(692) := std_logic_vector(to_signed(28609,16));
        tmp(693) := std_logic_vector(to_signed(28633,16));
        tmp(694) := std_logic_vector(to_signed(28658,16));
        tmp(695) := std_logic_vector(to_signed(28682,16));
        tmp(696) := std_logic_vector(to_signed(28706,16));
        tmp(697) := std_logic_vector(to_signed(28730,16));
        tmp(698) := std_logic_vector(to_signed(28755,16));
        tmp(699) := std_logic_vector(to_signed(28779,16));
        tmp(700) := std_logic_vector(to_signed(28803,16));
        tmp(701) := std_logic_vector(to_signed(28827,16));
        tmp(702) := std_logic_vector(to_signed(28850,16));
        tmp(703) := std_logic_vector(to_signed(28874,16));
        tmp(704) := std_logic_vector(to_signed(28898,16));
        tmp(705) := std_logic_vector(to_signed(28922,16));
        tmp(706) := std_logic_vector(to_signed(28945,16));
        tmp(707) := std_logic_vector(to_signed(28969,16));
        tmp(708) := std_logic_vector(to_signed(28992,16));
        tmp(709) := std_logic_vector(to_signed(29016,16));
        tmp(710) := std_logic_vector(to_signed(29039,16));
        tmp(711) := std_logic_vector(to_signed(29062,16));
        tmp(712) := std_logic_vector(to_signed(29085,16));
        tmp(713) := std_logic_vector(to_signed(29108,16));
        tmp(714) := std_logic_vector(to_signed(29131,16));
        tmp(715) := std_logic_vector(to_signed(29154,16));
        tmp(716) := std_logic_vector(to_signed(29177,16));
        tmp(717) := std_logic_vector(to_signed(29200,16));
        tmp(718) := std_logic_vector(to_signed(29223,16));
        tmp(719) := std_logic_vector(to_signed(29246,16));
        tmp(720) := std_logic_vector(to_signed(29268,16));
        tmp(721) := std_logic_vector(to_signed(29291,16));
        tmp(722) := std_logic_vector(to_signed(29313,16));
        tmp(723) := std_logic_vector(to_signed(29336,16));
        tmp(724) := std_logic_vector(to_signed(29358,16));
        tmp(725) := std_logic_vector(to_signed(29380,16));
        tmp(726) := std_logic_vector(to_signed(29403,16));
        tmp(727) := std_logic_vector(to_signed(29425,16));
        tmp(728) := std_logic_vector(to_signed(29447,16));
        tmp(729) := std_logic_vector(to_signed(29469,16));
        tmp(730) := std_logic_vector(to_signed(29491,16));
        tmp(731) := std_logic_vector(to_signed(29513,16));
        tmp(732) := std_logic_vector(to_signed(29534,16));
        tmp(733) := std_logic_vector(to_signed(29556,16));
        tmp(734) := std_logic_vector(to_signed(29578,16));
        tmp(735) := std_logic_vector(to_signed(29599,16));
        tmp(736) := std_logic_vector(to_signed(29621,16));
        tmp(737) := std_logic_vector(to_signed(29642,16));
        tmp(738) := std_logic_vector(to_signed(29664,16));
        tmp(739) := std_logic_vector(to_signed(29685,16));
        tmp(740) := std_logic_vector(to_signed(29706,16));
        tmp(741) := std_logic_vector(to_signed(29728,16));
        tmp(742) := std_logic_vector(to_signed(29749,16));
        tmp(743) := std_logic_vector(to_signed(29770,16));
        tmp(744) := std_logic_vector(to_signed(29791,16));
        tmp(745) := std_logic_vector(to_signed(29812,16));
        tmp(746) := std_logic_vector(to_signed(29832,16));
        tmp(747) := std_logic_vector(to_signed(29853,16));
        tmp(748) := std_logic_vector(to_signed(29874,16));
        tmp(749) := std_logic_vector(to_signed(29894,16));
        tmp(750) := std_logic_vector(to_signed(29915,16));
        tmp(751) := std_logic_vector(to_signed(29936,16));
        tmp(752) := std_logic_vector(to_signed(29956,16));
        tmp(753) := std_logic_vector(to_signed(29976,16));
        tmp(754) := std_logic_vector(to_signed(29997,16));
        tmp(755) := std_logic_vector(to_signed(30017,16));
        tmp(756) := std_logic_vector(to_signed(30037,16));
        tmp(757) := std_logic_vector(to_signed(30057,16));
        tmp(758) := std_logic_vector(to_signed(30077,16));
        tmp(759) := std_logic_vector(to_signed(30097,16));
        tmp(760) := std_logic_vector(to_signed(30117,16));
        tmp(761) := std_logic_vector(to_signed(30136,16));
        tmp(762) := std_logic_vector(to_signed(30156,16));
        tmp(763) := std_logic_vector(to_signed(30176,16));
        tmp(764) := std_logic_vector(to_signed(30195,16));
        tmp(765) := std_logic_vector(to_signed(30215,16));
        tmp(766) := std_logic_vector(to_signed(30234,16));
        tmp(767) := std_logic_vector(to_signed(30253,16));
        tmp(768) := std_logic_vector(to_signed(30273,16));
        tmp(769) := std_logic_vector(to_signed(30292,16));
        tmp(770) := std_logic_vector(to_signed(30311,16));
        tmp(771) := std_logic_vector(to_signed(30330,16));
        tmp(772) := std_logic_vector(to_signed(30349,16));
        tmp(773) := std_logic_vector(to_signed(30368,16));
        tmp(774) := std_logic_vector(to_signed(30387,16));
        tmp(775) := std_logic_vector(to_signed(30406,16));
        tmp(776) := std_logic_vector(to_signed(30424,16));
        tmp(777) := std_logic_vector(to_signed(30443,16));
        tmp(778) := std_logic_vector(to_signed(30462,16));
        tmp(779) := std_logic_vector(to_signed(30480,16));
        tmp(780) := std_logic_vector(to_signed(30498,16));
        tmp(781) := std_logic_vector(to_signed(30517,16));
        tmp(782) := std_logic_vector(to_signed(30535,16));
        tmp(783) := std_logic_vector(to_signed(30553,16));
        tmp(784) := std_logic_vector(to_signed(30571,16));
        tmp(785) := std_logic_vector(to_signed(30589,16));
        tmp(786) := std_logic_vector(to_signed(30607,16));
        tmp(787) := std_logic_vector(to_signed(30625,16));
        tmp(788) := std_logic_vector(to_signed(30643,16));
        tmp(789) := std_logic_vector(to_signed(30661,16));
        tmp(790) := std_logic_vector(to_signed(30679,16));
        tmp(791) := std_logic_vector(to_signed(30696,16));
        tmp(792) := std_logic_vector(to_signed(30714,16));
        tmp(793) := std_logic_vector(to_signed(30731,16));
        tmp(794) := std_logic_vector(to_signed(30749,16));
        tmp(795) := std_logic_vector(to_signed(30766,16));
        tmp(796) := std_logic_vector(to_signed(30783,16));
        tmp(797) := std_logic_vector(to_signed(30800,16));
        tmp(798) := std_logic_vector(to_signed(30818,16));
        tmp(799) := std_logic_vector(to_signed(30835,16));
        tmp(800) := std_logic_vector(to_signed(30852,16));
        tmp(801) := std_logic_vector(to_signed(30868,16));
        tmp(802) := std_logic_vector(to_signed(30885,16));
        tmp(803) := std_logic_vector(to_signed(30902,16));
        tmp(804) := std_logic_vector(to_signed(30919,16));
        tmp(805) := std_logic_vector(to_signed(30935,16));
        tmp(806) := std_logic_vector(to_signed(30952,16));
        tmp(807) := std_logic_vector(to_signed(30968,16));
        tmp(808) := std_logic_vector(to_signed(30985,16));
        tmp(809) := std_logic_vector(to_signed(31001,16));
        tmp(810) := std_logic_vector(to_signed(31017,16));
        tmp(811) := std_logic_vector(to_signed(31033,16));
        tmp(812) := std_logic_vector(to_signed(31050,16));
        tmp(813) := std_logic_vector(to_signed(31066,16));
        tmp(814) := std_logic_vector(to_signed(31082,16));
        tmp(815) := std_logic_vector(to_signed(31097,16));
        tmp(816) := std_logic_vector(to_signed(31113,16));
        tmp(817) := std_logic_vector(to_signed(31129,16));
        tmp(818) := std_logic_vector(to_signed(31145,16));
        tmp(819) := std_logic_vector(to_signed(31160,16));
        tmp(820) := std_logic_vector(to_signed(31176,16));
        tmp(821) := std_logic_vector(to_signed(31191,16));
        tmp(822) := std_logic_vector(to_signed(31206,16));
        tmp(823) := std_logic_vector(to_signed(31222,16));
        tmp(824) := std_logic_vector(to_signed(31237,16));
        tmp(825) := std_logic_vector(to_signed(31252,16));
        tmp(826) := std_logic_vector(to_signed(31267,16));
        tmp(827) := std_logic_vector(to_signed(31282,16));
        tmp(828) := std_logic_vector(to_signed(31297,16));
        tmp(829) := std_logic_vector(to_signed(31312,16));
        tmp(830) := std_logic_vector(to_signed(31327,16));
        tmp(831) := std_logic_vector(to_signed(31341,16));
        tmp(832) := std_logic_vector(to_signed(31356,16));
        tmp(833) := std_logic_vector(to_signed(31371,16));
        tmp(834) := std_logic_vector(to_signed(31385,16));
        tmp(835) := std_logic_vector(to_signed(31400,16));
        tmp(836) := std_logic_vector(to_signed(31414,16));
        tmp(837) := std_logic_vector(to_signed(31428,16));
        tmp(838) := std_logic_vector(to_signed(31442,16));
        tmp(839) := std_logic_vector(to_signed(31456,16));
        tmp(840) := std_logic_vector(to_signed(31470,16));
        tmp(841) := std_logic_vector(to_signed(31484,16));
        tmp(842) := std_logic_vector(to_signed(31498,16));
        tmp(843) := std_logic_vector(to_signed(31512,16));
        tmp(844) := std_logic_vector(to_signed(31526,16));
        tmp(845) := std_logic_vector(to_signed(31539,16));
        tmp(846) := std_logic_vector(to_signed(31553,16));
        tmp(847) := std_logic_vector(to_signed(31567,16));
        tmp(848) := std_logic_vector(to_signed(31580,16));
        tmp(849) := std_logic_vector(to_signed(31593,16));
        tmp(850) := std_logic_vector(to_signed(31607,16));
        tmp(851) := std_logic_vector(to_signed(31620,16));
        tmp(852) := std_logic_vector(to_signed(31633,16));
        tmp(853) := std_logic_vector(to_signed(31646,16));
        tmp(854) := std_logic_vector(to_signed(31659,16));
        tmp(855) := std_logic_vector(to_signed(31672,16));
        tmp(856) := std_logic_vector(to_signed(31685,16));
        tmp(857) := std_logic_vector(to_signed(31698,16));
        tmp(858) := std_logic_vector(to_signed(31710,16));
        tmp(859) := std_logic_vector(to_signed(31723,16));
        tmp(860) := std_logic_vector(to_signed(31736,16));
        tmp(861) := std_logic_vector(to_signed(31748,16));
        tmp(862) := std_logic_vector(to_signed(31760,16));
        tmp(863) := std_logic_vector(to_signed(31773,16));
        tmp(864) := std_logic_vector(to_signed(31785,16));
        tmp(865) := std_logic_vector(to_signed(31797,16));
        tmp(866) := std_logic_vector(to_signed(31809,16));
        tmp(867) := std_logic_vector(to_signed(31821,16));
        tmp(868) := std_logic_vector(to_signed(31833,16));
        tmp(869) := std_logic_vector(to_signed(31845,16));
        tmp(870) := std_logic_vector(to_signed(31857,16));
        tmp(871) := std_logic_vector(to_signed(31869,16));
        tmp(872) := std_logic_vector(to_signed(31880,16));
        tmp(873) := std_logic_vector(to_signed(31892,16));
        tmp(874) := std_logic_vector(to_signed(31903,16));
        tmp(875) := std_logic_vector(to_signed(31915,16));
        tmp(876) := std_logic_vector(to_signed(31926,16));
        tmp(877) := std_logic_vector(to_signed(31937,16));
        tmp(878) := std_logic_vector(to_signed(31949,16));
        tmp(879) := std_logic_vector(to_signed(31960,16));
        tmp(880) := std_logic_vector(to_signed(31971,16));
        tmp(881) := std_logic_vector(to_signed(31982,16));
        tmp(882) := std_logic_vector(to_signed(31993,16));
        tmp(883) := std_logic_vector(to_signed(32004,16));
        tmp(884) := std_logic_vector(to_signed(32014,16));
        tmp(885) := std_logic_vector(to_signed(32025,16));
        tmp(886) := std_logic_vector(to_signed(32036,16));
        tmp(887) := std_logic_vector(to_signed(32046,16));
        tmp(888) := std_logic_vector(to_signed(32057,16));
        tmp(889) := std_logic_vector(to_signed(32067,16));
        tmp(890) := std_logic_vector(to_signed(32077,16));
        tmp(891) := std_logic_vector(to_signed(32087,16));
        tmp(892) := std_logic_vector(to_signed(32098,16));
        tmp(893) := std_logic_vector(to_signed(32108,16));
        tmp(894) := std_logic_vector(to_signed(32118,16));
        tmp(895) := std_logic_vector(to_signed(32128,16));
        tmp(896) := std_logic_vector(to_signed(32137,16));
        tmp(897) := std_logic_vector(to_signed(32147,16));
        tmp(898) := std_logic_vector(to_signed(32157,16));
        tmp(899) := std_logic_vector(to_signed(32166,16));
        tmp(900) := std_logic_vector(to_signed(32176,16));
        tmp(901) := std_logic_vector(to_signed(32185,16));
        tmp(902) := std_logic_vector(to_signed(32195,16));
        tmp(903) := std_logic_vector(to_signed(32204,16));
        tmp(904) := std_logic_vector(to_signed(32213,16));
        tmp(905) := std_logic_vector(to_signed(32223,16));
        tmp(906) := std_logic_vector(to_signed(32232,16));
        tmp(907) := std_logic_vector(to_signed(32241,16));
        tmp(908) := std_logic_vector(to_signed(32250,16));
        tmp(909) := std_logic_vector(to_signed(32258,16));
        tmp(910) := std_logic_vector(to_signed(32267,16));
        tmp(911) := std_logic_vector(to_signed(32276,16));
        tmp(912) := std_logic_vector(to_signed(32285,16));
        tmp(913) := std_logic_vector(to_signed(32293,16));
        tmp(914) := std_logic_vector(to_signed(32302,16));
        tmp(915) := std_logic_vector(to_signed(32310,16));
        tmp(916) := std_logic_vector(to_signed(32318,16));
        tmp(917) := std_logic_vector(to_signed(32327,16));
        tmp(918) := std_logic_vector(to_signed(32335,16));
        tmp(919) := std_logic_vector(to_signed(32343,16));
        tmp(920) := std_logic_vector(to_signed(32351,16));
        tmp(921) := std_logic_vector(to_signed(32359,16));
        tmp(922) := std_logic_vector(to_signed(32367,16));
        tmp(923) := std_logic_vector(to_signed(32375,16));
        tmp(924) := std_logic_vector(to_signed(32382,16));
        tmp(925) := std_logic_vector(to_signed(32390,16));
        tmp(926) := std_logic_vector(to_signed(32397,16));
        tmp(927) := std_logic_vector(to_signed(32405,16));
        tmp(928) := std_logic_vector(to_signed(32412,16));
        tmp(929) := std_logic_vector(to_signed(32420,16));
        tmp(930) := std_logic_vector(to_signed(32427,16));
        tmp(931) := std_logic_vector(to_signed(32434,16));
        tmp(932) := std_logic_vector(to_signed(32441,16));
        tmp(933) := std_logic_vector(to_signed(32448,16));
        tmp(934) := std_logic_vector(to_signed(32455,16));
        tmp(935) := std_logic_vector(to_signed(32462,16));
        tmp(936) := std_logic_vector(to_signed(32469,16));
        tmp(937) := std_logic_vector(to_signed(32476,16));
        tmp(938) := std_logic_vector(to_signed(32482,16));
        tmp(939) := std_logic_vector(to_signed(32489,16));
        tmp(940) := std_logic_vector(to_signed(32495,16));
        tmp(941) := std_logic_vector(to_signed(32502,16));
        tmp(942) := std_logic_vector(to_signed(32508,16));
        tmp(943) := std_logic_vector(to_signed(32514,16));
        tmp(944) := std_logic_vector(to_signed(32521,16));
        tmp(945) := std_logic_vector(to_signed(32527,16));
        tmp(946) := std_logic_vector(to_signed(32533,16));
        tmp(947) := std_logic_vector(to_signed(32539,16));
        tmp(948) := std_logic_vector(to_signed(32545,16));
        tmp(949) := std_logic_vector(to_signed(32550,16));
        tmp(950) := std_logic_vector(to_signed(32556,16));
        tmp(951) := std_logic_vector(to_signed(32562,16));
        tmp(952) := std_logic_vector(to_signed(32567,16));
        tmp(953) := std_logic_vector(to_signed(32573,16));
        tmp(954) := std_logic_vector(to_signed(32578,16));
        tmp(955) := std_logic_vector(to_signed(32584,16));
        tmp(956) := std_logic_vector(to_signed(32589,16));
        tmp(957) := std_logic_vector(to_signed(32594,16));
        tmp(958) := std_logic_vector(to_signed(32599,16));
        tmp(959) := std_logic_vector(to_signed(32604,16));
        tmp(960) := std_logic_vector(to_signed(32609,16));
        tmp(961) := std_logic_vector(to_signed(32614,16));
        tmp(962) := std_logic_vector(to_signed(32619,16));
        tmp(963) := std_logic_vector(to_signed(32624,16));
        tmp(964) := std_logic_vector(to_signed(32628,16));
        tmp(965) := std_logic_vector(to_signed(32633,16));
        tmp(966) := std_logic_vector(to_signed(32637,16));
        tmp(967) := std_logic_vector(to_signed(32642,16));
        tmp(968) := std_logic_vector(to_signed(32646,16));
        tmp(969) := std_logic_vector(to_signed(32650,16));
        tmp(970) := std_logic_vector(to_signed(32655,16));
        tmp(971) := std_logic_vector(to_signed(32659,16));
        tmp(972) := std_logic_vector(to_signed(32663,16));
        tmp(973) := std_logic_vector(to_signed(32667,16));
        tmp(974) := std_logic_vector(to_signed(32671,16));
        tmp(975) := std_logic_vector(to_signed(32674,16));
        tmp(976) := std_logic_vector(to_signed(32678,16));
        tmp(977) := std_logic_vector(to_signed(32682,16));
        tmp(978) := std_logic_vector(to_signed(32685,16));
        tmp(979) := std_logic_vector(to_signed(32689,16));
        tmp(980) := std_logic_vector(to_signed(32692,16));
        tmp(981) := std_logic_vector(to_signed(32696,16));
        tmp(982) := std_logic_vector(to_signed(32699,16));
        tmp(983) := std_logic_vector(to_signed(32702,16));
        tmp(984) := std_logic_vector(to_signed(32705,16));
        tmp(985) := std_logic_vector(to_signed(32708,16));
        tmp(986) := std_logic_vector(to_signed(32711,16));
        tmp(987) := std_logic_vector(to_signed(32714,16));
        tmp(988) := std_logic_vector(to_signed(32717,16));
        tmp(989) := std_logic_vector(to_signed(32720,16));
        tmp(990) := std_logic_vector(to_signed(32722,16));
        tmp(991) := std_logic_vector(to_signed(32725,16));
        tmp(992) := std_logic_vector(to_signed(32728,16));
        tmp(993) := std_logic_vector(to_signed(32730,16));
        tmp(994) := std_logic_vector(to_signed(32732,16));
        tmp(995) := std_logic_vector(to_signed(32735,16));
        tmp(996) := std_logic_vector(to_signed(32737,16));
        tmp(997) := std_logic_vector(to_signed(32739,16));
        tmp(998) := std_logic_vector(to_signed(32741,16));
        tmp(999) := std_logic_vector(to_signed(32743,16));
        tmp(1000) := std_logic_vector(to_signed(32745,16));
        tmp(1001) := std_logic_vector(to_signed(32747,16));
        tmp(1002) := std_logic_vector(to_signed(32748,16));
        tmp(1003) := std_logic_vector(to_signed(32750,16));
        tmp(1004) := std_logic_vector(to_signed(32752,16));
        tmp(1005) := std_logic_vector(to_signed(32753,16));
        tmp(1006) := std_logic_vector(to_signed(32755,16));
        tmp(1007) := std_logic_vector(to_signed(32756,16));
        tmp(1008) := std_logic_vector(to_signed(32757,16));
        tmp(1009) := std_logic_vector(to_signed(32758,16));
        tmp(1010) := std_logic_vector(to_signed(32759,16));
        tmp(1011) := std_logic_vector(to_signed(32760,16));
        tmp(1012) := std_logic_vector(to_signed(32761,16));
        tmp(1013) := std_logic_vector(to_signed(32762,16));
        tmp(1014) := std_logic_vector(to_signed(32763,16));
        tmp(1015) := std_logic_vector(to_signed(32764,16));
        tmp(1016) := std_logic_vector(to_signed(32765,16));
        tmp(1017) := std_logic_vector(to_signed(32765,16));
        tmp(1018) := std_logic_vector(to_signed(32766,16));
        tmp(1019) := std_logic_vector(to_signed(32766,16));
        tmp(1020) := std_logic_vector(to_signed(32766,16));
        tmp(1021) := std_logic_vector(to_signed(32767,16));
        tmp(1022) := std_logic_vector(to_signed(32767,16));
        tmp(1023) := std_logic_vector(to_signed(32767,16));
        tmp(1024) := std_logic_vector(to_signed(32767,16));
        tmp(1025) := std_logic_vector(to_signed(32767,16));
        tmp(1026) := std_logic_vector(to_signed(32767,16));
        tmp(1027) := std_logic_vector(to_signed(32767,16));
        tmp(1028) := std_logic_vector(to_signed(32766,16));
        tmp(1029) := std_logic_vector(to_signed(32766,16));
        tmp(1030) := std_logic_vector(to_signed(32766,16));
        tmp(1031) := std_logic_vector(to_signed(32765,16));
        tmp(1032) := std_logic_vector(to_signed(32765,16));
        tmp(1033) := std_logic_vector(to_signed(32764,16));
        tmp(1034) := std_logic_vector(to_signed(32763,16));
        tmp(1035) := std_logic_vector(to_signed(32762,16));
        tmp(1036) := std_logic_vector(to_signed(32761,16));
        tmp(1037) := std_logic_vector(to_signed(32760,16));
        tmp(1038) := std_logic_vector(to_signed(32759,16));
        tmp(1039) := std_logic_vector(to_signed(32758,16));
        tmp(1040) := std_logic_vector(to_signed(32757,16));
        tmp(1041) := std_logic_vector(to_signed(32756,16));
        tmp(1042) := std_logic_vector(to_signed(32755,16));
        tmp(1043) := std_logic_vector(to_signed(32753,16));
        tmp(1044) := std_logic_vector(to_signed(32752,16));
        tmp(1045) := std_logic_vector(to_signed(32750,16));
        tmp(1046) := std_logic_vector(to_signed(32748,16));
        tmp(1047) := std_logic_vector(to_signed(32747,16));
        tmp(1048) := std_logic_vector(to_signed(32745,16));
        tmp(1049) := std_logic_vector(to_signed(32743,16));
        tmp(1050) := std_logic_vector(to_signed(32741,16));
        tmp(1051) := std_logic_vector(to_signed(32739,16));
        tmp(1052) := std_logic_vector(to_signed(32737,16));
        tmp(1053) := std_logic_vector(to_signed(32735,16));
        tmp(1054) := std_logic_vector(to_signed(32732,16));
        tmp(1055) := std_logic_vector(to_signed(32730,16));
        tmp(1056) := std_logic_vector(to_signed(32728,16));
        tmp(1057) := std_logic_vector(to_signed(32725,16));
        tmp(1058) := std_logic_vector(to_signed(32722,16));
        tmp(1059) := std_logic_vector(to_signed(32720,16));
        tmp(1060) := std_logic_vector(to_signed(32717,16));
        tmp(1061) := std_logic_vector(to_signed(32714,16));
        tmp(1062) := std_logic_vector(to_signed(32711,16));
        tmp(1063) := std_logic_vector(to_signed(32708,16));
        tmp(1064) := std_logic_vector(to_signed(32705,16));
        tmp(1065) := std_logic_vector(to_signed(32702,16));
        tmp(1066) := std_logic_vector(to_signed(32699,16));
        tmp(1067) := std_logic_vector(to_signed(32696,16));
        tmp(1068) := std_logic_vector(to_signed(32692,16));
        tmp(1069) := std_logic_vector(to_signed(32689,16));
        tmp(1070) := std_logic_vector(to_signed(32685,16));
        tmp(1071) := std_logic_vector(to_signed(32682,16));
        tmp(1072) := std_logic_vector(to_signed(32678,16));
        tmp(1073) := std_logic_vector(to_signed(32674,16));
        tmp(1074) := std_logic_vector(to_signed(32671,16));
        tmp(1075) := std_logic_vector(to_signed(32667,16));
        tmp(1076) := std_logic_vector(to_signed(32663,16));
        tmp(1077) := std_logic_vector(to_signed(32659,16));
        tmp(1078) := std_logic_vector(to_signed(32655,16));
        tmp(1079) := std_logic_vector(to_signed(32650,16));
        tmp(1080) := std_logic_vector(to_signed(32646,16));
        tmp(1081) := std_logic_vector(to_signed(32642,16));
        tmp(1082) := std_logic_vector(to_signed(32637,16));
        tmp(1083) := std_logic_vector(to_signed(32633,16));
        tmp(1084) := std_logic_vector(to_signed(32628,16));
        tmp(1085) := std_logic_vector(to_signed(32624,16));
        tmp(1086) := std_logic_vector(to_signed(32619,16));
        tmp(1087) := std_logic_vector(to_signed(32614,16));
        tmp(1088) := std_logic_vector(to_signed(32609,16));
        tmp(1089) := std_logic_vector(to_signed(32604,16));
        tmp(1090) := std_logic_vector(to_signed(32599,16));
        tmp(1091) := std_logic_vector(to_signed(32594,16));
        tmp(1092) := std_logic_vector(to_signed(32589,16));
        tmp(1093) := std_logic_vector(to_signed(32584,16));
        tmp(1094) := std_logic_vector(to_signed(32578,16));
        tmp(1095) := std_logic_vector(to_signed(32573,16));
        tmp(1096) := std_logic_vector(to_signed(32567,16));
        tmp(1097) := std_logic_vector(to_signed(32562,16));
        tmp(1098) := std_logic_vector(to_signed(32556,16));
        tmp(1099) := std_logic_vector(to_signed(32550,16));
        tmp(1100) := std_logic_vector(to_signed(32545,16));
        tmp(1101) := std_logic_vector(to_signed(32539,16));
        tmp(1102) := std_logic_vector(to_signed(32533,16));
        tmp(1103) := std_logic_vector(to_signed(32527,16));
        tmp(1104) := std_logic_vector(to_signed(32521,16));
        tmp(1105) := std_logic_vector(to_signed(32514,16));
        tmp(1106) := std_logic_vector(to_signed(32508,16));
        tmp(1107) := std_logic_vector(to_signed(32502,16));
        tmp(1108) := std_logic_vector(to_signed(32495,16));
        tmp(1109) := std_logic_vector(to_signed(32489,16));
        tmp(1110) := std_logic_vector(to_signed(32482,16));
        tmp(1111) := std_logic_vector(to_signed(32476,16));
        tmp(1112) := std_logic_vector(to_signed(32469,16));
        tmp(1113) := std_logic_vector(to_signed(32462,16));
        tmp(1114) := std_logic_vector(to_signed(32455,16));
        tmp(1115) := std_logic_vector(to_signed(32448,16));
        tmp(1116) := std_logic_vector(to_signed(32441,16));
        tmp(1117) := std_logic_vector(to_signed(32434,16));
        tmp(1118) := std_logic_vector(to_signed(32427,16));
        tmp(1119) := std_logic_vector(to_signed(32420,16));
        tmp(1120) := std_logic_vector(to_signed(32412,16));
        tmp(1121) := std_logic_vector(to_signed(32405,16));
        tmp(1122) := std_logic_vector(to_signed(32397,16));
        tmp(1123) := std_logic_vector(to_signed(32390,16));
        tmp(1124) := std_logic_vector(to_signed(32382,16));
        tmp(1125) := std_logic_vector(to_signed(32375,16));
        tmp(1126) := std_logic_vector(to_signed(32367,16));
        tmp(1127) := std_logic_vector(to_signed(32359,16));
        tmp(1128) := std_logic_vector(to_signed(32351,16));
        tmp(1129) := std_logic_vector(to_signed(32343,16));
        tmp(1130) := std_logic_vector(to_signed(32335,16));
        tmp(1131) := std_logic_vector(to_signed(32327,16));
        tmp(1132) := std_logic_vector(to_signed(32318,16));
        tmp(1133) := std_logic_vector(to_signed(32310,16));
        tmp(1134) := std_logic_vector(to_signed(32302,16));
        tmp(1135) := std_logic_vector(to_signed(32293,16));
        tmp(1136) := std_logic_vector(to_signed(32285,16));
        tmp(1137) := std_logic_vector(to_signed(32276,16));
        tmp(1138) := std_logic_vector(to_signed(32267,16));
        tmp(1139) := std_logic_vector(to_signed(32258,16));
        tmp(1140) := std_logic_vector(to_signed(32250,16));
        tmp(1141) := std_logic_vector(to_signed(32241,16));
        tmp(1142) := std_logic_vector(to_signed(32232,16));
        tmp(1143) := std_logic_vector(to_signed(32223,16));
        tmp(1144) := std_logic_vector(to_signed(32213,16));
        tmp(1145) := std_logic_vector(to_signed(32204,16));
        tmp(1146) := std_logic_vector(to_signed(32195,16));
        tmp(1147) := std_logic_vector(to_signed(32185,16));
        tmp(1148) := std_logic_vector(to_signed(32176,16));
        tmp(1149) := std_logic_vector(to_signed(32166,16));
        tmp(1150) := std_logic_vector(to_signed(32157,16));
        tmp(1151) := std_logic_vector(to_signed(32147,16));
        tmp(1152) := std_logic_vector(to_signed(32137,16));
        tmp(1153) := std_logic_vector(to_signed(32128,16));
        tmp(1154) := std_logic_vector(to_signed(32118,16));
        tmp(1155) := std_logic_vector(to_signed(32108,16));
        tmp(1156) := std_logic_vector(to_signed(32098,16));
        tmp(1157) := std_logic_vector(to_signed(32087,16));
        tmp(1158) := std_logic_vector(to_signed(32077,16));
        tmp(1159) := std_logic_vector(to_signed(32067,16));
        tmp(1160) := std_logic_vector(to_signed(32057,16));
        tmp(1161) := std_logic_vector(to_signed(32046,16));
        tmp(1162) := std_logic_vector(to_signed(32036,16));
        tmp(1163) := std_logic_vector(to_signed(32025,16));
        tmp(1164) := std_logic_vector(to_signed(32014,16));
        tmp(1165) := std_logic_vector(to_signed(32004,16));
        tmp(1166) := std_logic_vector(to_signed(31993,16));
        tmp(1167) := std_logic_vector(to_signed(31982,16));
        tmp(1168) := std_logic_vector(to_signed(31971,16));
        tmp(1169) := std_logic_vector(to_signed(31960,16));
        tmp(1170) := std_logic_vector(to_signed(31949,16));
        tmp(1171) := std_logic_vector(to_signed(31937,16));
        tmp(1172) := std_logic_vector(to_signed(31926,16));
        tmp(1173) := std_logic_vector(to_signed(31915,16));
        tmp(1174) := std_logic_vector(to_signed(31903,16));
        tmp(1175) := std_logic_vector(to_signed(31892,16));
        tmp(1176) := std_logic_vector(to_signed(31880,16));
        tmp(1177) := std_logic_vector(to_signed(31869,16));
        tmp(1178) := std_logic_vector(to_signed(31857,16));
        tmp(1179) := std_logic_vector(to_signed(31845,16));
        tmp(1180) := std_logic_vector(to_signed(31833,16));
        tmp(1181) := std_logic_vector(to_signed(31821,16));
        tmp(1182) := std_logic_vector(to_signed(31809,16));
        tmp(1183) := std_logic_vector(to_signed(31797,16));
        tmp(1184) := std_logic_vector(to_signed(31785,16));
        tmp(1185) := std_logic_vector(to_signed(31773,16));
        tmp(1186) := std_logic_vector(to_signed(31760,16));
        tmp(1187) := std_logic_vector(to_signed(31748,16));
        tmp(1188) := std_logic_vector(to_signed(31736,16));
        tmp(1189) := std_logic_vector(to_signed(31723,16));
        tmp(1190) := std_logic_vector(to_signed(31710,16));
        tmp(1191) := std_logic_vector(to_signed(31698,16));
        tmp(1192) := std_logic_vector(to_signed(31685,16));
        tmp(1193) := std_logic_vector(to_signed(31672,16));
        tmp(1194) := std_logic_vector(to_signed(31659,16));
        tmp(1195) := std_logic_vector(to_signed(31646,16));
        tmp(1196) := std_logic_vector(to_signed(31633,16));
        tmp(1197) := std_logic_vector(to_signed(31620,16));
        tmp(1198) := std_logic_vector(to_signed(31607,16));
        tmp(1199) := std_logic_vector(to_signed(31593,16));
        tmp(1200) := std_logic_vector(to_signed(31580,16));
        tmp(1201) := std_logic_vector(to_signed(31567,16));
        tmp(1202) := std_logic_vector(to_signed(31553,16));
        tmp(1203) := std_logic_vector(to_signed(31539,16));
        tmp(1204) := std_logic_vector(to_signed(31526,16));
        tmp(1205) := std_logic_vector(to_signed(31512,16));
        tmp(1206) := std_logic_vector(to_signed(31498,16));
        tmp(1207) := std_logic_vector(to_signed(31484,16));
        tmp(1208) := std_logic_vector(to_signed(31470,16));
        tmp(1209) := std_logic_vector(to_signed(31456,16));
        tmp(1210) := std_logic_vector(to_signed(31442,16));
        tmp(1211) := std_logic_vector(to_signed(31428,16));
        tmp(1212) := std_logic_vector(to_signed(31414,16));
        tmp(1213) := std_logic_vector(to_signed(31400,16));
        tmp(1214) := std_logic_vector(to_signed(31385,16));
        tmp(1215) := std_logic_vector(to_signed(31371,16));
        tmp(1216) := std_logic_vector(to_signed(31356,16));
        tmp(1217) := std_logic_vector(to_signed(31341,16));
        tmp(1218) := std_logic_vector(to_signed(31327,16));
        tmp(1219) := std_logic_vector(to_signed(31312,16));
        tmp(1220) := std_logic_vector(to_signed(31297,16));
        tmp(1221) := std_logic_vector(to_signed(31282,16));
        tmp(1222) := std_logic_vector(to_signed(31267,16));
        tmp(1223) := std_logic_vector(to_signed(31252,16));
        tmp(1224) := std_logic_vector(to_signed(31237,16));
        tmp(1225) := std_logic_vector(to_signed(31222,16));
        tmp(1226) := std_logic_vector(to_signed(31206,16));
        tmp(1227) := std_logic_vector(to_signed(31191,16));
        tmp(1228) := std_logic_vector(to_signed(31176,16));
        tmp(1229) := std_logic_vector(to_signed(31160,16));
        tmp(1230) := std_logic_vector(to_signed(31145,16));
        tmp(1231) := std_logic_vector(to_signed(31129,16));
        tmp(1232) := std_logic_vector(to_signed(31113,16));
        tmp(1233) := std_logic_vector(to_signed(31097,16));
        tmp(1234) := std_logic_vector(to_signed(31082,16));
        tmp(1235) := std_logic_vector(to_signed(31066,16));
        tmp(1236) := std_logic_vector(to_signed(31050,16));
        tmp(1237) := std_logic_vector(to_signed(31033,16));
        tmp(1238) := std_logic_vector(to_signed(31017,16));
        tmp(1239) := std_logic_vector(to_signed(31001,16));
        tmp(1240) := std_logic_vector(to_signed(30985,16));
        tmp(1241) := std_logic_vector(to_signed(30968,16));
        tmp(1242) := std_logic_vector(to_signed(30952,16));
        tmp(1243) := std_logic_vector(to_signed(30935,16));
        tmp(1244) := std_logic_vector(to_signed(30919,16));
        tmp(1245) := std_logic_vector(to_signed(30902,16));
        tmp(1246) := std_logic_vector(to_signed(30885,16));
        tmp(1247) := std_logic_vector(to_signed(30868,16));
        tmp(1248) := std_logic_vector(to_signed(30852,16));
        tmp(1249) := std_logic_vector(to_signed(30835,16));
        tmp(1250) := std_logic_vector(to_signed(30818,16));
        tmp(1251) := std_logic_vector(to_signed(30800,16));
        tmp(1252) := std_logic_vector(to_signed(30783,16));
        tmp(1253) := std_logic_vector(to_signed(30766,16));
        tmp(1254) := std_logic_vector(to_signed(30749,16));
        tmp(1255) := std_logic_vector(to_signed(30731,16));
        tmp(1256) := std_logic_vector(to_signed(30714,16));
        tmp(1257) := std_logic_vector(to_signed(30696,16));
        tmp(1258) := std_logic_vector(to_signed(30679,16));
        tmp(1259) := std_logic_vector(to_signed(30661,16));
        tmp(1260) := std_logic_vector(to_signed(30643,16));
        tmp(1261) := std_logic_vector(to_signed(30625,16));
        tmp(1262) := std_logic_vector(to_signed(30607,16));
        tmp(1263) := std_logic_vector(to_signed(30589,16));
        tmp(1264) := std_logic_vector(to_signed(30571,16));
        tmp(1265) := std_logic_vector(to_signed(30553,16));
        tmp(1266) := std_logic_vector(to_signed(30535,16));
        tmp(1267) := std_logic_vector(to_signed(30517,16));
        tmp(1268) := std_logic_vector(to_signed(30498,16));
        tmp(1269) := std_logic_vector(to_signed(30480,16));
        tmp(1270) := std_logic_vector(to_signed(30462,16));
        tmp(1271) := std_logic_vector(to_signed(30443,16));
        tmp(1272) := std_logic_vector(to_signed(30424,16));
        tmp(1273) := std_logic_vector(to_signed(30406,16));
        tmp(1274) := std_logic_vector(to_signed(30387,16));
        tmp(1275) := std_logic_vector(to_signed(30368,16));
        tmp(1276) := std_logic_vector(to_signed(30349,16));
        tmp(1277) := std_logic_vector(to_signed(30330,16));
        tmp(1278) := std_logic_vector(to_signed(30311,16));
        tmp(1279) := std_logic_vector(to_signed(30292,16));
        tmp(1280) := std_logic_vector(to_signed(30273,16));
        tmp(1281) := std_logic_vector(to_signed(30253,16));
        tmp(1282) := std_logic_vector(to_signed(30234,16));
        tmp(1283) := std_logic_vector(to_signed(30215,16));
        tmp(1284) := std_logic_vector(to_signed(30195,16));
        tmp(1285) := std_logic_vector(to_signed(30176,16));
        tmp(1286) := std_logic_vector(to_signed(30156,16));
        tmp(1287) := std_logic_vector(to_signed(30136,16));
        tmp(1288) := std_logic_vector(to_signed(30117,16));
        tmp(1289) := std_logic_vector(to_signed(30097,16));
        tmp(1290) := std_logic_vector(to_signed(30077,16));
        tmp(1291) := std_logic_vector(to_signed(30057,16));
        tmp(1292) := std_logic_vector(to_signed(30037,16));
        tmp(1293) := std_logic_vector(to_signed(30017,16));
        tmp(1294) := std_logic_vector(to_signed(29997,16));
        tmp(1295) := std_logic_vector(to_signed(29976,16));
        tmp(1296) := std_logic_vector(to_signed(29956,16));
        tmp(1297) := std_logic_vector(to_signed(29936,16));
        tmp(1298) := std_logic_vector(to_signed(29915,16));
        tmp(1299) := std_logic_vector(to_signed(29894,16));
        tmp(1300) := std_logic_vector(to_signed(29874,16));
        tmp(1301) := std_logic_vector(to_signed(29853,16));
        tmp(1302) := std_logic_vector(to_signed(29832,16));
        tmp(1303) := std_logic_vector(to_signed(29812,16));
        tmp(1304) := std_logic_vector(to_signed(29791,16));
        tmp(1305) := std_logic_vector(to_signed(29770,16));
        tmp(1306) := std_logic_vector(to_signed(29749,16));
        tmp(1307) := std_logic_vector(to_signed(29728,16));
        tmp(1308) := std_logic_vector(to_signed(29706,16));
        tmp(1309) := std_logic_vector(to_signed(29685,16));
        tmp(1310) := std_logic_vector(to_signed(29664,16));
        tmp(1311) := std_logic_vector(to_signed(29642,16));
        tmp(1312) := std_logic_vector(to_signed(29621,16));
        tmp(1313) := std_logic_vector(to_signed(29599,16));
        tmp(1314) := std_logic_vector(to_signed(29578,16));
        tmp(1315) := std_logic_vector(to_signed(29556,16));
        tmp(1316) := std_logic_vector(to_signed(29534,16));
        tmp(1317) := std_logic_vector(to_signed(29513,16));
        tmp(1318) := std_logic_vector(to_signed(29491,16));
        tmp(1319) := std_logic_vector(to_signed(29469,16));
        tmp(1320) := std_logic_vector(to_signed(29447,16));
        tmp(1321) := std_logic_vector(to_signed(29425,16));
        tmp(1322) := std_logic_vector(to_signed(29403,16));
        tmp(1323) := std_logic_vector(to_signed(29380,16));
        tmp(1324) := std_logic_vector(to_signed(29358,16));
        tmp(1325) := std_logic_vector(to_signed(29336,16));
        tmp(1326) := std_logic_vector(to_signed(29313,16));
        tmp(1327) := std_logic_vector(to_signed(29291,16));
        tmp(1328) := std_logic_vector(to_signed(29268,16));
        tmp(1329) := std_logic_vector(to_signed(29246,16));
        tmp(1330) := std_logic_vector(to_signed(29223,16));
        tmp(1331) := std_logic_vector(to_signed(29200,16));
        tmp(1332) := std_logic_vector(to_signed(29177,16));
        tmp(1333) := std_logic_vector(to_signed(29154,16));
        tmp(1334) := std_logic_vector(to_signed(29131,16));
        tmp(1335) := std_logic_vector(to_signed(29108,16));
        tmp(1336) := std_logic_vector(to_signed(29085,16));
        tmp(1337) := std_logic_vector(to_signed(29062,16));
        tmp(1338) := std_logic_vector(to_signed(29039,16));
        tmp(1339) := std_logic_vector(to_signed(29016,16));
        tmp(1340) := std_logic_vector(to_signed(28992,16));
        tmp(1341) := std_logic_vector(to_signed(28969,16));
        tmp(1342) := std_logic_vector(to_signed(28945,16));
        tmp(1343) := std_logic_vector(to_signed(28922,16));
        tmp(1344) := std_logic_vector(to_signed(28898,16));
        tmp(1345) := std_logic_vector(to_signed(28874,16));
        tmp(1346) := std_logic_vector(to_signed(28850,16));
        tmp(1347) := std_logic_vector(to_signed(28827,16));
        tmp(1348) := std_logic_vector(to_signed(28803,16));
        tmp(1349) := std_logic_vector(to_signed(28779,16));
        tmp(1350) := std_logic_vector(to_signed(28755,16));
        tmp(1351) := std_logic_vector(to_signed(28730,16));
        tmp(1352) := std_logic_vector(to_signed(28706,16));
        tmp(1353) := std_logic_vector(to_signed(28682,16));
        tmp(1354) := std_logic_vector(to_signed(28658,16));
        tmp(1355) := std_logic_vector(to_signed(28633,16));
        tmp(1356) := std_logic_vector(to_signed(28609,16));
        tmp(1357) := std_logic_vector(to_signed(28584,16));
        tmp(1358) := std_logic_vector(to_signed(28560,16));
        tmp(1359) := std_logic_vector(to_signed(28535,16));
        tmp(1360) := std_logic_vector(to_signed(28510,16));
        tmp(1361) := std_logic_vector(to_signed(28485,16));
        tmp(1362) := std_logic_vector(to_signed(28460,16));
        tmp(1363) := std_logic_vector(to_signed(28436,16));
        tmp(1364) := std_logic_vector(to_signed(28411,16));
        tmp(1365) := std_logic_vector(to_signed(28385,16));
        tmp(1366) := std_logic_vector(to_signed(28360,16));
        tmp(1367) := std_logic_vector(to_signed(28335,16));
        tmp(1368) := std_logic_vector(to_signed(28310,16));
        tmp(1369) := std_logic_vector(to_signed(28284,16));
        tmp(1370) := std_logic_vector(to_signed(28259,16));
        tmp(1371) := std_logic_vector(to_signed(28234,16));
        tmp(1372) := std_logic_vector(to_signed(28208,16));
        tmp(1373) := std_logic_vector(to_signed(28182,16));
        tmp(1374) := std_logic_vector(to_signed(28157,16));
        tmp(1375) := std_logic_vector(to_signed(28131,16));
        tmp(1376) := std_logic_vector(to_signed(28105,16));
        tmp(1377) := std_logic_vector(to_signed(28079,16));
        tmp(1378) := std_logic_vector(to_signed(28053,16));
        tmp(1379) := std_logic_vector(to_signed(28027,16));
        tmp(1380) := std_logic_vector(to_signed(28001,16));
        tmp(1381) := std_logic_vector(to_signed(27975,16));
        tmp(1382) := std_logic_vector(to_signed(27949,16));
        tmp(1383) := std_logic_vector(to_signed(27923,16));
        tmp(1384) := std_logic_vector(to_signed(27896,16));
        tmp(1385) := std_logic_vector(to_signed(27870,16));
        tmp(1386) := std_logic_vector(to_signed(27843,16));
        tmp(1387) := std_logic_vector(to_signed(27817,16));
        tmp(1388) := std_logic_vector(to_signed(27790,16));
        tmp(1389) := std_logic_vector(to_signed(27764,16));
        tmp(1390) := std_logic_vector(to_signed(27737,16));
        tmp(1391) := std_logic_vector(to_signed(27710,16));
        tmp(1392) := std_logic_vector(to_signed(27683,16));
        tmp(1393) := std_logic_vector(to_signed(27656,16));
        tmp(1394) := std_logic_vector(to_signed(27629,16));
        tmp(1395) := std_logic_vector(to_signed(27602,16));
        tmp(1396) := std_logic_vector(to_signed(27575,16));
        tmp(1397) := std_logic_vector(to_signed(27548,16));
        tmp(1398) := std_logic_vector(to_signed(27521,16));
        tmp(1399) := std_logic_vector(to_signed(27493,16));
        tmp(1400) := std_logic_vector(to_signed(27466,16));
        tmp(1401) := std_logic_vector(to_signed(27439,16));
        tmp(1402) := std_logic_vector(to_signed(27411,16));
        tmp(1403) := std_logic_vector(to_signed(27384,16));
        tmp(1404) := std_logic_vector(to_signed(27356,16));
        tmp(1405) := std_logic_vector(to_signed(27328,16));
        tmp(1406) := std_logic_vector(to_signed(27300,16));
        tmp(1407) := std_logic_vector(to_signed(27273,16));
        tmp(1408) := std_logic_vector(to_signed(27245,16));
        tmp(1409) := std_logic_vector(to_signed(27217,16));
        tmp(1410) := std_logic_vector(to_signed(27189,16));
        tmp(1411) := std_logic_vector(to_signed(27161,16));
        tmp(1412) := std_logic_vector(to_signed(27133,16));
        tmp(1413) := std_logic_vector(to_signed(27104,16));
        tmp(1414) := std_logic_vector(to_signed(27076,16));
        tmp(1415) := std_logic_vector(to_signed(27048,16));
        tmp(1416) := std_logic_vector(to_signed(27019,16));
        tmp(1417) := std_logic_vector(to_signed(26991,16));
        tmp(1418) := std_logic_vector(to_signed(26962,16));
        tmp(1419) := std_logic_vector(to_signed(26934,16));
        tmp(1420) := std_logic_vector(to_signed(26905,16));
        tmp(1421) := std_logic_vector(to_signed(26876,16));
        tmp(1422) := std_logic_vector(to_signed(26848,16));
        tmp(1423) := std_logic_vector(to_signed(26819,16));
        tmp(1424) := std_logic_vector(to_signed(26790,16));
        tmp(1425) := std_logic_vector(to_signed(26761,16));
        tmp(1426) := std_logic_vector(to_signed(26732,16));
        tmp(1427) := std_logic_vector(to_signed(26703,16));
        tmp(1428) := std_logic_vector(to_signed(26674,16));
        tmp(1429) := std_logic_vector(to_signed(26644,16));
        tmp(1430) := std_logic_vector(to_signed(26615,16));
        tmp(1431) := std_logic_vector(to_signed(26586,16));
        tmp(1432) := std_logic_vector(to_signed(26556,16));
        tmp(1433) := std_logic_vector(to_signed(26527,16));
        tmp(1434) := std_logic_vector(to_signed(26497,16));
        tmp(1435) := std_logic_vector(to_signed(26468,16));
        tmp(1436) := std_logic_vector(to_signed(26438,16));
        tmp(1437) := std_logic_vector(to_signed(26408,16));
        tmp(1438) := std_logic_vector(to_signed(26378,16));
        tmp(1439) := std_logic_vector(to_signed(26349,16));
        tmp(1440) := std_logic_vector(to_signed(26319,16));
        tmp(1441) := std_logic_vector(to_signed(26289,16));
        tmp(1442) := std_logic_vector(to_signed(26259,16));
        tmp(1443) := std_logic_vector(to_signed(26229,16));
        tmp(1444) := std_logic_vector(to_signed(26198,16));
        tmp(1445) := std_logic_vector(to_signed(26168,16));
        tmp(1446) := std_logic_vector(to_signed(26138,16));
        tmp(1447) := std_logic_vector(to_signed(26108,16));
        tmp(1448) := std_logic_vector(to_signed(26077,16));
        tmp(1449) := std_logic_vector(to_signed(26047,16));
        tmp(1450) := std_logic_vector(to_signed(26016,16));
        tmp(1451) := std_logic_vector(to_signed(25986,16));
        tmp(1452) := std_logic_vector(to_signed(25955,16));
        tmp(1453) := std_logic_vector(to_signed(25924,16));
        tmp(1454) := std_logic_vector(to_signed(25893,16));
        tmp(1455) := std_logic_vector(to_signed(25863,16));
        tmp(1456) := std_logic_vector(to_signed(25832,16));
        tmp(1457) := std_logic_vector(to_signed(25801,16));
        tmp(1458) := std_logic_vector(to_signed(25770,16));
        tmp(1459) := std_logic_vector(to_signed(25739,16));
        tmp(1460) := std_logic_vector(to_signed(25708,16));
        tmp(1461) := std_logic_vector(to_signed(25676,16));
        tmp(1462) := std_logic_vector(to_signed(25645,16));
        tmp(1463) := std_logic_vector(to_signed(25614,16));
        tmp(1464) := std_logic_vector(to_signed(25582,16));
        tmp(1465) := std_logic_vector(to_signed(25551,16));
        tmp(1466) := std_logic_vector(to_signed(25519,16));
        tmp(1467) := std_logic_vector(to_signed(25488,16));
        tmp(1468) := std_logic_vector(to_signed(25456,16));
        tmp(1469) := std_logic_vector(to_signed(25425,16));
        tmp(1470) := std_logic_vector(to_signed(25393,16));
        tmp(1471) := std_logic_vector(to_signed(25361,16));
        tmp(1472) := std_logic_vector(to_signed(25329,16));
        tmp(1473) := std_logic_vector(to_signed(25297,16));
        tmp(1474) := std_logic_vector(to_signed(25265,16));
        tmp(1475) := std_logic_vector(to_signed(25233,16));
        tmp(1476) := std_logic_vector(to_signed(25201,16));
        tmp(1477) := std_logic_vector(to_signed(25169,16));
        tmp(1478) := std_logic_vector(to_signed(25137,16));
        tmp(1479) := std_logic_vector(to_signed(25105,16));
        tmp(1480) := std_logic_vector(to_signed(25072,16));
        tmp(1481) := std_logic_vector(to_signed(25040,16));
        tmp(1482) := std_logic_vector(to_signed(25007,16));
        tmp(1483) := std_logic_vector(to_signed(24975,16));
        tmp(1484) := std_logic_vector(to_signed(24942,16));
        tmp(1485) := std_logic_vector(to_signed(24910,16));
        tmp(1486) := std_logic_vector(to_signed(24877,16));
        tmp(1487) := std_logic_vector(to_signed(24844,16));
        tmp(1488) := std_logic_vector(to_signed(24811,16));
        tmp(1489) := std_logic_vector(to_signed(24779,16));
        tmp(1490) := std_logic_vector(to_signed(24746,16));
        tmp(1491) := std_logic_vector(to_signed(24713,16));
        tmp(1492) := std_logic_vector(to_signed(24680,16));
        tmp(1493) := std_logic_vector(to_signed(24647,16));
        tmp(1494) := std_logic_vector(to_signed(24613,16));
        tmp(1495) := std_logic_vector(to_signed(24580,16));
        tmp(1496) := std_logic_vector(to_signed(24547,16));
        tmp(1497) := std_logic_vector(to_signed(24514,16));
        tmp(1498) := std_logic_vector(to_signed(24480,16));
        tmp(1499) := std_logic_vector(to_signed(24447,16));
        tmp(1500) := std_logic_vector(to_signed(24413,16));
        tmp(1501) := std_logic_vector(to_signed(24380,16));
        tmp(1502) := std_logic_vector(to_signed(24346,16));
        tmp(1503) := std_logic_vector(to_signed(24312,16));
        tmp(1504) := std_logic_vector(to_signed(24279,16));
        tmp(1505) := std_logic_vector(to_signed(24245,16));
        tmp(1506) := std_logic_vector(to_signed(24211,16));
        tmp(1507) := std_logic_vector(to_signed(24177,16));
        tmp(1508) := std_logic_vector(to_signed(24143,16));
        tmp(1509) := std_logic_vector(to_signed(24109,16));
        tmp(1510) := std_logic_vector(to_signed(24075,16));
        tmp(1511) := std_logic_vector(to_signed(24041,16));
        tmp(1512) := std_logic_vector(to_signed(24007,16));
        tmp(1513) := std_logic_vector(to_signed(23973,16));
        tmp(1514) := std_logic_vector(to_signed(23938,16));
        tmp(1515) := std_logic_vector(to_signed(23904,16));
        tmp(1516) := std_logic_vector(to_signed(23870,16));
        tmp(1517) := std_logic_vector(to_signed(23835,16));
        tmp(1518) := std_logic_vector(to_signed(23801,16));
        tmp(1519) := std_logic_vector(to_signed(23766,16));
        tmp(1520) := std_logic_vector(to_signed(23731,16));
        tmp(1521) := std_logic_vector(to_signed(23697,16));
        tmp(1522) := std_logic_vector(to_signed(23662,16));
        tmp(1523) := std_logic_vector(to_signed(23627,16));
        tmp(1524) := std_logic_vector(to_signed(23592,16));
        tmp(1525) := std_logic_vector(to_signed(23557,16));
        tmp(1526) := std_logic_vector(to_signed(23522,16));
        tmp(1527) := std_logic_vector(to_signed(23487,16));
        tmp(1528) := std_logic_vector(to_signed(23452,16));
        tmp(1529) := std_logic_vector(to_signed(23417,16));
        tmp(1530) := std_logic_vector(to_signed(23382,16));
        tmp(1531) := std_logic_vector(to_signed(23347,16));
        tmp(1532) := std_logic_vector(to_signed(23311,16));
        tmp(1533) := std_logic_vector(to_signed(23276,16));
        tmp(1534) := std_logic_vector(to_signed(23241,16));
        tmp(1535) := std_logic_vector(to_signed(23205,16));
        tmp(1536) := std_logic_vector(to_signed(23170,16));
        tmp(1537) := std_logic_vector(to_signed(23134,16));
        tmp(1538) := std_logic_vector(to_signed(23099,16));
        tmp(1539) := std_logic_vector(to_signed(23063,16));
        tmp(1540) := std_logic_vector(to_signed(23027,16));
        tmp(1541) := std_logic_vector(to_signed(22991,16));
        tmp(1542) := std_logic_vector(to_signed(22956,16));
        tmp(1543) := std_logic_vector(to_signed(22920,16));
        tmp(1544) := std_logic_vector(to_signed(22884,16));
        tmp(1545) := std_logic_vector(to_signed(22848,16));
        tmp(1546) := std_logic_vector(to_signed(22812,16));
        tmp(1547) := std_logic_vector(to_signed(22776,16));
        tmp(1548) := std_logic_vector(to_signed(22739,16));
        tmp(1549) := std_logic_vector(to_signed(22703,16));
        tmp(1550) := std_logic_vector(to_signed(22667,16));
        tmp(1551) := std_logic_vector(to_signed(22631,16));
        tmp(1552) := std_logic_vector(to_signed(22594,16));
        tmp(1553) := std_logic_vector(to_signed(22558,16));
        tmp(1554) := std_logic_vector(to_signed(22521,16));
        tmp(1555) := std_logic_vector(to_signed(22485,16));
        tmp(1556) := std_logic_vector(to_signed(22448,16));
        tmp(1557) := std_logic_vector(to_signed(22411,16));
        tmp(1558) := std_logic_vector(to_signed(22375,16));
        tmp(1559) := std_logic_vector(to_signed(22338,16));
        tmp(1560) := std_logic_vector(to_signed(22301,16));
        tmp(1561) := std_logic_vector(to_signed(22264,16));
        tmp(1562) := std_logic_vector(to_signed(22227,16));
        tmp(1563) := std_logic_vector(to_signed(22191,16));
        tmp(1564) := std_logic_vector(to_signed(22154,16));
        tmp(1565) := std_logic_vector(to_signed(22116,16));
        tmp(1566) := std_logic_vector(to_signed(22079,16));
        tmp(1567) := std_logic_vector(to_signed(22042,16));
        tmp(1568) := std_logic_vector(to_signed(22005,16));
        tmp(1569) := std_logic_vector(to_signed(21968,16));
        tmp(1570) := std_logic_vector(to_signed(21930,16));
        tmp(1571) := std_logic_vector(to_signed(21893,16));
        tmp(1572) := std_logic_vector(to_signed(21856,16));
        tmp(1573) := std_logic_vector(to_signed(21818,16));
        tmp(1574) := std_logic_vector(to_signed(21781,16));
        tmp(1575) := std_logic_vector(to_signed(21743,16));
        tmp(1576) := std_logic_vector(to_signed(21705,16));
        tmp(1577) := std_logic_vector(to_signed(21668,16));
        tmp(1578) := std_logic_vector(to_signed(21630,16));
        tmp(1579) := std_logic_vector(to_signed(21592,16));
        tmp(1580) := std_logic_vector(to_signed(21554,16));
        tmp(1581) := std_logic_vector(to_signed(21516,16));
        tmp(1582) := std_logic_vector(to_signed(21479,16));
        tmp(1583) := std_logic_vector(to_signed(21441,16));
        tmp(1584) := std_logic_vector(to_signed(21403,16));
        tmp(1585) := std_logic_vector(to_signed(21364,16));
        tmp(1586) := std_logic_vector(to_signed(21326,16));
        tmp(1587) := std_logic_vector(to_signed(21288,16));
        tmp(1588) := std_logic_vector(to_signed(21250,16));
        tmp(1589) := std_logic_vector(to_signed(21212,16));
        tmp(1590) := std_logic_vector(to_signed(21173,16));
        tmp(1591) := std_logic_vector(to_signed(21135,16));
        tmp(1592) := std_logic_vector(to_signed(21096,16));
        tmp(1593) := std_logic_vector(to_signed(21058,16));
        tmp(1594) := std_logic_vector(to_signed(21019,16));
        tmp(1595) := std_logic_vector(to_signed(20981,16));
        tmp(1596) := std_logic_vector(to_signed(20942,16));
        tmp(1597) := std_logic_vector(to_signed(20904,16));
        tmp(1598) := std_logic_vector(to_signed(20865,16));
        tmp(1599) := std_logic_vector(to_signed(20826,16));
        tmp(1600) := std_logic_vector(to_signed(20787,16));
        tmp(1601) := std_logic_vector(to_signed(20748,16));
        tmp(1602) := std_logic_vector(to_signed(20709,16));
        tmp(1603) := std_logic_vector(to_signed(20670,16));
        tmp(1604) := std_logic_vector(to_signed(20631,16));
        tmp(1605) := std_logic_vector(to_signed(20592,16));
        tmp(1606) := std_logic_vector(to_signed(20553,16));
        tmp(1607) := std_logic_vector(to_signed(20514,16));
        tmp(1608) := std_logic_vector(to_signed(20475,16));
        tmp(1609) := std_logic_vector(to_signed(20436,16));
        tmp(1610) := std_logic_vector(to_signed(20396,16));
        tmp(1611) := std_logic_vector(to_signed(20357,16));
        tmp(1612) := std_logic_vector(to_signed(20317,16));
        tmp(1613) := std_logic_vector(to_signed(20278,16));
        tmp(1614) := std_logic_vector(to_signed(20238,16));
        tmp(1615) := std_logic_vector(to_signed(20199,16));
        tmp(1616) := std_logic_vector(to_signed(20159,16));
        tmp(1617) := std_logic_vector(to_signed(20120,16));
        tmp(1618) := std_logic_vector(to_signed(20080,16));
        tmp(1619) := std_logic_vector(to_signed(20040,16));
        tmp(1620) := std_logic_vector(to_signed(20000,16));
        tmp(1621) := std_logic_vector(to_signed(19961,16));
        tmp(1622) := std_logic_vector(to_signed(19921,16));
        tmp(1623) := std_logic_vector(to_signed(19881,16));
        tmp(1624) := std_logic_vector(to_signed(19841,16));
        tmp(1625) := std_logic_vector(to_signed(19801,16));
        tmp(1626) := std_logic_vector(to_signed(19761,16));
        tmp(1627) := std_logic_vector(to_signed(19721,16));
        tmp(1628) := std_logic_vector(to_signed(19680,16));
        tmp(1629) := std_logic_vector(to_signed(19640,16));
        tmp(1630) := std_logic_vector(to_signed(19600,16));
        tmp(1631) := std_logic_vector(to_signed(19560,16));
        tmp(1632) := std_logic_vector(to_signed(19519,16));
        tmp(1633) := std_logic_vector(to_signed(19479,16));
        tmp(1634) := std_logic_vector(to_signed(19438,16));
        tmp(1635) := std_logic_vector(to_signed(19398,16));
        tmp(1636) := std_logic_vector(to_signed(19357,16));
        tmp(1637) := std_logic_vector(to_signed(19317,16));
        tmp(1638) := std_logic_vector(to_signed(19276,16));
        tmp(1639) := std_logic_vector(to_signed(19236,16));
        tmp(1640) := std_logic_vector(to_signed(19195,16));
        tmp(1641) := std_logic_vector(to_signed(19154,16));
        tmp(1642) := std_logic_vector(to_signed(19113,16));
        tmp(1643) := std_logic_vector(to_signed(19072,16));
        tmp(1644) := std_logic_vector(to_signed(19032,16));
        tmp(1645) := std_logic_vector(to_signed(18991,16));
        tmp(1646) := std_logic_vector(to_signed(18950,16));
        tmp(1647) := std_logic_vector(to_signed(18909,16));
        tmp(1648) := std_logic_vector(to_signed(18868,16));
        tmp(1649) := std_logic_vector(to_signed(18826,16));
        tmp(1650) := std_logic_vector(to_signed(18785,16));
        tmp(1651) := std_logic_vector(to_signed(18744,16));
        tmp(1652) := std_logic_vector(to_signed(18703,16));
        tmp(1653) := std_logic_vector(to_signed(18661,16));
        tmp(1654) := std_logic_vector(to_signed(18620,16));
        tmp(1655) := std_logic_vector(to_signed(18579,16));
        tmp(1656) := std_logic_vector(to_signed(18537,16));
        tmp(1657) := std_logic_vector(to_signed(18496,16));
        tmp(1658) := std_logic_vector(to_signed(18454,16));
        tmp(1659) := std_logic_vector(to_signed(18413,16));
        tmp(1660) := std_logic_vector(to_signed(18371,16));
        tmp(1661) := std_logic_vector(to_signed(18330,16));
        tmp(1662) := std_logic_vector(to_signed(18288,16));
        tmp(1663) := std_logic_vector(to_signed(18246,16));
        tmp(1664) := std_logic_vector(to_signed(18204,16));
        tmp(1665) := std_logic_vector(to_signed(18163,16));
        tmp(1666) := std_logic_vector(to_signed(18121,16));
        tmp(1667) := std_logic_vector(to_signed(18079,16));
        tmp(1668) := std_logic_vector(to_signed(18037,16));
        tmp(1669) := std_logic_vector(to_signed(17995,16));
        tmp(1670) := std_logic_vector(to_signed(17953,16));
        tmp(1671) := std_logic_vector(to_signed(17911,16));
        tmp(1672) := std_logic_vector(to_signed(17869,16));
        tmp(1673) := std_logic_vector(to_signed(17827,16));
        tmp(1674) := std_logic_vector(to_signed(17784,16));
        tmp(1675) := std_logic_vector(to_signed(17742,16));
        tmp(1676) := std_logic_vector(to_signed(17700,16));
        tmp(1677) := std_logic_vector(to_signed(17657,16));
        tmp(1678) := std_logic_vector(to_signed(17615,16));
        tmp(1679) := std_logic_vector(to_signed(17573,16));
        tmp(1680) := std_logic_vector(to_signed(17530,16));
        tmp(1681) := std_logic_vector(to_signed(17488,16));
        tmp(1682) := std_logic_vector(to_signed(17445,16));
        tmp(1683) := std_logic_vector(to_signed(17403,16));
        tmp(1684) := std_logic_vector(to_signed(17360,16));
        tmp(1685) := std_logic_vector(to_signed(17317,16));
        tmp(1686) := std_logic_vector(to_signed(17275,16));
        tmp(1687) := std_logic_vector(to_signed(17232,16));
        tmp(1688) := std_logic_vector(to_signed(17189,16));
        tmp(1689) := std_logic_vector(to_signed(17146,16));
        tmp(1690) := std_logic_vector(to_signed(17104,16));
        tmp(1691) := std_logic_vector(to_signed(17061,16));
        tmp(1692) := std_logic_vector(to_signed(17018,16));
        tmp(1693) := std_logic_vector(to_signed(16975,16));
        tmp(1694) := std_logic_vector(to_signed(16932,16));
        tmp(1695) := std_logic_vector(to_signed(16889,16));
        tmp(1696) := std_logic_vector(to_signed(16846,16));
        tmp(1697) := std_logic_vector(to_signed(16802,16));
        tmp(1698) := std_logic_vector(to_signed(16759,16));
        tmp(1699) := std_logic_vector(to_signed(16716,16));
        tmp(1700) := std_logic_vector(to_signed(16673,16));
        tmp(1701) := std_logic_vector(to_signed(16630,16));
        tmp(1702) := std_logic_vector(to_signed(16586,16));
        tmp(1703) := std_logic_vector(to_signed(16543,16));
        tmp(1704) := std_logic_vector(to_signed(16499,16));
        tmp(1705) := std_logic_vector(to_signed(16456,16));
        tmp(1706) := std_logic_vector(to_signed(16413,16));
        tmp(1707) := std_logic_vector(to_signed(16369,16));
        tmp(1708) := std_logic_vector(to_signed(16325,16));
        tmp(1709) := std_logic_vector(to_signed(16282,16));
        tmp(1710) := std_logic_vector(to_signed(16238,16));
        tmp(1711) := std_logic_vector(to_signed(16195,16));
        tmp(1712) := std_logic_vector(to_signed(16151,16));
        tmp(1713) := std_logic_vector(to_signed(16107,16));
        tmp(1714) := std_logic_vector(to_signed(16063,16));
        tmp(1715) := std_logic_vector(to_signed(16019,16));
        tmp(1716) := std_logic_vector(to_signed(15976,16));
        tmp(1717) := std_logic_vector(to_signed(15932,16));
        tmp(1718) := std_logic_vector(to_signed(15888,16));
        tmp(1719) := std_logic_vector(to_signed(15844,16));
        tmp(1720) := std_logic_vector(to_signed(15800,16));
        tmp(1721) := std_logic_vector(to_signed(15756,16));
        tmp(1722) := std_logic_vector(to_signed(15712,16));
        tmp(1723) := std_logic_vector(to_signed(15667,16));
        tmp(1724) := std_logic_vector(to_signed(15623,16));
        tmp(1725) := std_logic_vector(to_signed(15579,16));
        tmp(1726) := std_logic_vector(to_signed(15535,16));
        tmp(1727) := std_logic_vector(to_signed(15491,16));
        tmp(1728) := std_logic_vector(to_signed(15446,16));
        tmp(1729) := std_logic_vector(to_signed(15402,16));
        tmp(1730) := std_logic_vector(to_signed(15358,16));
        tmp(1731) := std_logic_vector(to_signed(15313,16));
        tmp(1732) := std_logic_vector(to_signed(15269,16));
        tmp(1733) := std_logic_vector(to_signed(15224,16));
        tmp(1734) := std_logic_vector(to_signed(15180,16));
        tmp(1735) := std_logic_vector(to_signed(15135,16));
        tmp(1736) := std_logic_vector(to_signed(15090,16));
        tmp(1737) := std_logic_vector(to_signed(15046,16));
        tmp(1738) := std_logic_vector(to_signed(15001,16));
        tmp(1739) := std_logic_vector(to_signed(14956,16));
        tmp(1740) := std_logic_vector(to_signed(14912,16));
        tmp(1741) := std_logic_vector(to_signed(14867,16));
        tmp(1742) := std_logic_vector(to_signed(14822,16));
        tmp(1743) := std_logic_vector(to_signed(14777,16));
        tmp(1744) := std_logic_vector(to_signed(14732,16));
        tmp(1745) := std_logic_vector(to_signed(14688,16));
        tmp(1746) := std_logic_vector(to_signed(14643,16));
        tmp(1747) := std_logic_vector(to_signed(14598,16));
        tmp(1748) := std_logic_vector(to_signed(14553,16));
        tmp(1749) := std_logic_vector(to_signed(14507,16));
        tmp(1750) := std_logic_vector(to_signed(14462,16));
        tmp(1751) := std_logic_vector(to_signed(14417,16));
        tmp(1752) := std_logic_vector(to_signed(14372,16));
        tmp(1753) := std_logic_vector(to_signed(14327,16));
        tmp(1754) := std_logic_vector(to_signed(14282,16));
        tmp(1755) := std_logic_vector(to_signed(14236,16));
        tmp(1756) := std_logic_vector(to_signed(14191,16));
        tmp(1757) := std_logic_vector(to_signed(14146,16));
        tmp(1758) := std_logic_vector(to_signed(14101,16));
        tmp(1759) := std_logic_vector(to_signed(14055,16));
        tmp(1760) := std_logic_vector(to_signed(14010,16));
        tmp(1761) := std_logic_vector(to_signed(13964,16));
        tmp(1762) := std_logic_vector(to_signed(13919,16));
        tmp(1763) := std_logic_vector(to_signed(13873,16));
        tmp(1764) := std_logic_vector(to_signed(13828,16));
        tmp(1765) := std_logic_vector(to_signed(13782,16));
        tmp(1766) := std_logic_vector(to_signed(13736,16));
        tmp(1767) := std_logic_vector(to_signed(13691,16));
        tmp(1768) := std_logic_vector(to_signed(13645,16));
        tmp(1769) := std_logic_vector(to_signed(13599,16));
        tmp(1770) := std_logic_vector(to_signed(13554,16));
        tmp(1771) := std_logic_vector(to_signed(13508,16));
        tmp(1772) := std_logic_vector(to_signed(13462,16));
        tmp(1773) := std_logic_vector(to_signed(13416,16));
        tmp(1774) := std_logic_vector(to_signed(13370,16));
        tmp(1775) := std_logic_vector(to_signed(13324,16));
        tmp(1776) := std_logic_vector(to_signed(13279,16));
        tmp(1777) := std_logic_vector(to_signed(13233,16));
        tmp(1778) := std_logic_vector(to_signed(13187,16));
        tmp(1779) := std_logic_vector(to_signed(13141,16));
        tmp(1780) := std_logic_vector(to_signed(13094,16));
        tmp(1781) := std_logic_vector(to_signed(13048,16));
        tmp(1782) := std_logic_vector(to_signed(13002,16));
        tmp(1783) := std_logic_vector(to_signed(12956,16));
        tmp(1784) := std_logic_vector(to_signed(12910,16));
        tmp(1785) := std_logic_vector(to_signed(12864,16));
        tmp(1786) := std_logic_vector(to_signed(12817,16));
        tmp(1787) := std_logic_vector(to_signed(12771,16));
        tmp(1788) := std_logic_vector(to_signed(12725,16));
        tmp(1789) := std_logic_vector(to_signed(12679,16));
        tmp(1790) := std_logic_vector(to_signed(12632,16));
        tmp(1791) := std_logic_vector(to_signed(12586,16));
        tmp(1792) := std_logic_vector(to_signed(12539,16));
        tmp(1793) := std_logic_vector(to_signed(12493,16));
        tmp(1794) := std_logic_vector(to_signed(12446,16));
        tmp(1795) := std_logic_vector(to_signed(12400,16));
        tmp(1796) := std_logic_vector(to_signed(12353,16));
        tmp(1797) := std_logic_vector(to_signed(12307,16));
        tmp(1798) := std_logic_vector(to_signed(12260,16));
        tmp(1799) := std_logic_vector(to_signed(12214,16));
        tmp(1800) := std_logic_vector(to_signed(12167,16));
        tmp(1801) := std_logic_vector(to_signed(12120,16));
        tmp(1802) := std_logic_vector(to_signed(12074,16));
        tmp(1803) := std_logic_vector(to_signed(12027,16));
        tmp(1804) := std_logic_vector(to_signed(11980,16));
        tmp(1805) := std_logic_vector(to_signed(11933,16));
        tmp(1806) := std_logic_vector(to_signed(11886,16));
        tmp(1807) := std_logic_vector(to_signed(11840,16));
        tmp(1808) := std_logic_vector(to_signed(11793,16));
        tmp(1809) := std_logic_vector(to_signed(11746,16));
        tmp(1810) := std_logic_vector(to_signed(11699,16));
        tmp(1811) := std_logic_vector(to_signed(11652,16));
        tmp(1812) := std_logic_vector(to_signed(11605,16));
        tmp(1813) := std_logic_vector(to_signed(11558,16));
        tmp(1814) := std_logic_vector(to_signed(11511,16));
        tmp(1815) := std_logic_vector(to_signed(11464,16));
        tmp(1816) := std_logic_vector(to_signed(11417,16));
        tmp(1817) := std_logic_vector(to_signed(11370,16));
        tmp(1818) := std_logic_vector(to_signed(11322,16));
        tmp(1819) := std_logic_vector(to_signed(11275,16));
        tmp(1820) := std_logic_vector(to_signed(11228,16));
        tmp(1821) := std_logic_vector(to_signed(11181,16));
        tmp(1822) := std_logic_vector(to_signed(11133,16));
        tmp(1823) := std_logic_vector(to_signed(11086,16));
        tmp(1824) := std_logic_vector(to_signed(11039,16));
        tmp(1825) := std_logic_vector(to_signed(10992,16));
        tmp(1826) := std_logic_vector(to_signed(10944,16));
        tmp(1827) := std_logic_vector(to_signed(10897,16));
        tmp(1828) := std_logic_vector(to_signed(10849,16));
        tmp(1829) := std_logic_vector(to_signed(10802,16));
        tmp(1830) := std_logic_vector(to_signed(10754,16));
        tmp(1831) := std_logic_vector(to_signed(10707,16));
        tmp(1832) := std_logic_vector(to_signed(10659,16));
        tmp(1833) := std_logic_vector(to_signed(10612,16));
        tmp(1834) := std_logic_vector(to_signed(10564,16));
        tmp(1835) := std_logic_vector(to_signed(10517,16));
        tmp(1836) := std_logic_vector(to_signed(10469,16));
        tmp(1837) := std_logic_vector(to_signed(10421,16));
        tmp(1838) := std_logic_vector(to_signed(10374,16));
        tmp(1839) := std_logic_vector(to_signed(10326,16));
        tmp(1840) := std_logic_vector(to_signed(10278,16));
        tmp(1841) := std_logic_vector(to_signed(10231,16));
        tmp(1842) := std_logic_vector(to_signed(10183,16));
        tmp(1843) := std_logic_vector(to_signed(10135,16));
        tmp(1844) := std_logic_vector(to_signed(10087,16));
        tmp(1845) := std_logic_vector(to_signed(10039,16));
        tmp(1846) := std_logic_vector(to_signed(9992,16));
        tmp(1847) := std_logic_vector(to_signed(9944,16));
        tmp(1848) := std_logic_vector(to_signed(9896,16));
        tmp(1849) := std_logic_vector(to_signed(9848,16));
        tmp(1850) := std_logic_vector(to_signed(9800,16));
        tmp(1851) := std_logic_vector(to_signed(9752,16));
        tmp(1852) := std_logic_vector(to_signed(9704,16));
        tmp(1853) := std_logic_vector(to_signed(9656,16));
        tmp(1854) := std_logic_vector(to_signed(9608,16));
        tmp(1855) := std_logic_vector(to_signed(9560,16));
        tmp(1856) := std_logic_vector(to_signed(9512,16));
        tmp(1857) := std_logic_vector(to_signed(9464,16));
        tmp(1858) := std_logic_vector(to_signed(9416,16));
        tmp(1859) := std_logic_vector(to_signed(9367,16));
        tmp(1860) := std_logic_vector(to_signed(9319,16));
        tmp(1861) := std_logic_vector(to_signed(9271,16));
        tmp(1862) := std_logic_vector(to_signed(9223,16));
        tmp(1863) := std_logic_vector(to_signed(9175,16));
        tmp(1864) := std_logic_vector(to_signed(9126,16));
        tmp(1865) := std_logic_vector(to_signed(9078,16));
        tmp(1866) := std_logic_vector(to_signed(9030,16));
        tmp(1867) := std_logic_vector(to_signed(8981,16));
        tmp(1868) := std_logic_vector(to_signed(8933,16));
        tmp(1869) := std_logic_vector(to_signed(8885,16));
        tmp(1870) := std_logic_vector(to_signed(8836,16));
        tmp(1871) := std_logic_vector(to_signed(8788,16));
        tmp(1872) := std_logic_vector(to_signed(8739,16));
        tmp(1873) := std_logic_vector(to_signed(8691,16));
        tmp(1874) := std_logic_vector(to_signed(8642,16));
        tmp(1875) := std_logic_vector(to_signed(8594,16));
        tmp(1876) := std_logic_vector(to_signed(8545,16));
        tmp(1877) := std_logic_vector(to_signed(8497,16));
        tmp(1878) := std_logic_vector(to_signed(8448,16));
        tmp(1879) := std_logic_vector(to_signed(8400,16));
        tmp(1880) := std_logic_vector(to_signed(8351,16));
        tmp(1881) := std_logic_vector(to_signed(8303,16));
        tmp(1882) := std_logic_vector(to_signed(8254,16));
        tmp(1883) := std_logic_vector(to_signed(8205,16));
        tmp(1884) := std_logic_vector(to_signed(8157,16));
        tmp(1885) := std_logic_vector(to_signed(8108,16));
        tmp(1886) := std_logic_vector(to_signed(8059,16));
        tmp(1887) := std_logic_vector(to_signed(8010,16));
        tmp(1888) := std_logic_vector(to_signed(7962,16));
        tmp(1889) := std_logic_vector(to_signed(7913,16));
        tmp(1890) := std_logic_vector(to_signed(7864,16));
        tmp(1891) := std_logic_vector(to_signed(7815,16));
        tmp(1892) := std_logic_vector(to_signed(7767,16));
        tmp(1893) := std_logic_vector(to_signed(7718,16));
        tmp(1894) := std_logic_vector(to_signed(7669,16));
        tmp(1895) := std_logic_vector(to_signed(7620,16));
        tmp(1896) := std_logic_vector(to_signed(7571,16));
        tmp(1897) := std_logic_vector(to_signed(7522,16));
        tmp(1898) := std_logic_vector(to_signed(7473,16));
        tmp(1899) := std_logic_vector(to_signed(7424,16));
        tmp(1900) := std_logic_vector(to_signed(7375,16));
        tmp(1901) := std_logic_vector(to_signed(7326,16));
        tmp(1902) := std_logic_vector(to_signed(7277,16));
        tmp(1903) := std_logic_vector(to_signed(7228,16));
        tmp(1904) := std_logic_vector(to_signed(7179,16));
        tmp(1905) := std_logic_vector(to_signed(7130,16));
        tmp(1906) := std_logic_vector(to_signed(7081,16));
        tmp(1907) := std_logic_vector(to_signed(7032,16));
        tmp(1908) := std_logic_vector(to_signed(6983,16));
        tmp(1909) := std_logic_vector(to_signed(6934,16));
        tmp(1910) := std_logic_vector(to_signed(6885,16));
        tmp(1911) := std_logic_vector(to_signed(6836,16));
        tmp(1912) := std_logic_vector(to_signed(6786,16));
        tmp(1913) := std_logic_vector(to_signed(6737,16));
        tmp(1914) := std_logic_vector(to_signed(6688,16));
        tmp(1915) := std_logic_vector(to_signed(6639,16));
        tmp(1916) := std_logic_vector(to_signed(6590,16));
        tmp(1917) := std_logic_vector(to_signed(6540,16));
        tmp(1918) := std_logic_vector(to_signed(6491,16));
        tmp(1919) := std_logic_vector(to_signed(6442,16));
        tmp(1920) := std_logic_vector(to_signed(6393,16));
        tmp(1921) := std_logic_vector(to_signed(6343,16));
        tmp(1922) := std_logic_vector(to_signed(6294,16));
        tmp(1923) := std_logic_vector(to_signed(6245,16));
        tmp(1924) := std_logic_vector(to_signed(6195,16));
        tmp(1925) := std_logic_vector(to_signed(6146,16));
        tmp(1926) := std_logic_vector(to_signed(6096,16));
        tmp(1927) := std_logic_vector(to_signed(6047,16));
        tmp(1928) := std_logic_vector(to_signed(5998,16));
        tmp(1929) := std_logic_vector(to_signed(5948,16));
        tmp(1930) := std_logic_vector(to_signed(5899,16));
        tmp(1931) := std_logic_vector(to_signed(5849,16));
        tmp(1932) := std_logic_vector(to_signed(5800,16));
        tmp(1933) := std_logic_vector(to_signed(5750,16));
        tmp(1934) := std_logic_vector(to_signed(5701,16));
        tmp(1935) := std_logic_vector(to_signed(5651,16));
        tmp(1936) := std_logic_vector(to_signed(5602,16));
        tmp(1937) := std_logic_vector(to_signed(5552,16));
        tmp(1938) := std_logic_vector(to_signed(5503,16));
        tmp(1939) := std_logic_vector(to_signed(5453,16));
        tmp(1940) := std_logic_vector(to_signed(5404,16));
        tmp(1941) := std_logic_vector(to_signed(5354,16));
        tmp(1942) := std_logic_vector(to_signed(5305,16));
        tmp(1943) := std_logic_vector(to_signed(5255,16));
        tmp(1944) := std_logic_vector(to_signed(5205,16));
        tmp(1945) := std_logic_vector(to_signed(5156,16));
        tmp(1946) := std_logic_vector(to_signed(5106,16));
        tmp(1947) := std_logic_vector(to_signed(5056,16));
        tmp(1948) := std_logic_vector(to_signed(5007,16));
        tmp(1949) := std_logic_vector(to_signed(4957,16));
        tmp(1950) := std_logic_vector(to_signed(4907,16));
        tmp(1951) := std_logic_vector(to_signed(4858,16));
        tmp(1952) := std_logic_vector(to_signed(4808,16));
        tmp(1953) := std_logic_vector(to_signed(4758,16));
        tmp(1954) := std_logic_vector(to_signed(4708,16));
        tmp(1955) := std_logic_vector(to_signed(4659,16));
        tmp(1956) := std_logic_vector(to_signed(4609,16));
        tmp(1957) := std_logic_vector(to_signed(4559,16));
        tmp(1958) := std_logic_vector(to_signed(4509,16));
        tmp(1959) := std_logic_vector(to_signed(4460,16));
        tmp(1960) := std_logic_vector(to_signed(4410,16));
        tmp(1961) := std_logic_vector(to_signed(4360,16));
        tmp(1962) := std_logic_vector(to_signed(4310,16));
        tmp(1963) := std_logic_vector(to_signed(4260,16));
        tmp(1964) := std_logic_vector(to_signed(4210,16));
        tmp(1965) := std_logic_vector(to_signed(4161,16));
        tmp(1966) := std_logic_vector(to_signed(4111,16));
        tmp(1967) := std_logic_vector(to_signed(4061,16));
        tmp(1968) := std_logic_vector(to_signed(4011,16));
        tmp(1969) := std_logic_vector(to_signed(3961,16));
        tmp(1970) := std_logic_vector(to_signed(3911,16));
        tmp(1971) := std_logic_vector(to_signed(3861,16));
        tmp(1972) := std_logic_vector(to_signed(3811,16));
        tmp(1973) := std_logic_vector(to_signed(3761,16));
        tmp(1974) := std_logic_vector(to_signed(3712,16));
        tmp(1975) := std_logic_vector(to_signed(3662,16));
        tmp(1976) := std_logic_vector(to_signed(3612,16));
        tmp(1977) := std_logic_vector(to_signed(3562,16));
        tmp(1978) := std_logic_vector(to_signed(3512,16));
        tmp(1979) := std_logic_vector(to_signed(3462,16));
        tmp(1980) := std_logic_vector(to_signed(3412,16));
        tmp(1981) := std_logic_vector(to_signed(3362,16));
        tmp(1982) := std_logic_vector(to_signed(3312,16));
        tmp(1983) := std_logic_vector(to_signed(3262,16));
        tmp(1984) := std_logic_vector(to_signed(3212,16));
        tmp(1985) := std_logic_vector(to_signed(3162,16));
        tmp(1986) := std_logic_vector(to_signed(3112,16));
        tmp(1987) := std_logic_vector(to_signed(3062,16));
        tmp(1988) := std_logic_vector(to_signed(3012,16));
        tmp(1989) := std_logic_vector(to_signed(2962,16));
        tmp(1990) := std_logic_vector(to_signed(2911,16));
        tmp(1991) := std_logic_vector(to_signed(2861,16));
        tmp(1992) := std_logic_vector(to_signed(2811,16));
        tmp(1993) := std_logic_vector(to_signed(2761,16));
        tmp(1994) := std_logic_vector(to_signed(2711,16));
        tmp(1995) := std_logic_vector(to_signed(2661,16));
        tmp(1996) := std_logic_vector(to_signed(2611,16));
        tmp(1997) := std_logic_vector(to_signed(2561,16));
        tmp(1998) := std_logic_vector(to_signed(2511,16));
        tmp(1999) := std_logic_vector(to_signed(2461,16));
        tmp(2000) := std_logic_vector(to_signed(2410,16));
        tmp(2001) := std_logic_vector(to_signed(2360,16));
        tmp(2002) := std_logic_vector(to_signed(2310,16));
        tmp(2003) := std_logic_vector(to_signed(2260,16));
        tmp(2004) := std_logic_vector(to_signed(2210,16));
        tmp(2005) := std_logic_vector(to_signed(2160,16));
        tmp(2006) := std_logic_vector(to_signed(2110,16));
        tmp(2007) := std_logic_vector(to_signed(2059,16));
        tmp(2008) := std_logic_vector(to_signed(2009,16));
        tmp(2009) := std_logic_vector(to_signed(1959,16));
        tmp(2010) := std_logic_vector(to_signed(1909,16));
        tmp(2011) := std_logic_vector(to_signed(1859,16));
        tmp(2012) := std_logic_vector(to_signed(1809,16));
        tmp(2013) := std_logic_vector(to_signed(1758,16));
        tmp(2014) := std_logic_vector(to_signed(1708,16));
        tmp(2015) := std_logic_vector(to_signed(1658,16));
        tmp(2016) := std_logic_vector(to_signed(1608,16));
        tmp(2017) := std_logic_vector(to_signed(1558,16));
        tmp(2018) := std_logic_vector(to_signed(1507,16));
        tmp(2019) := std_logic_vector(to_signed(1457,16));
        tmp(2020) := std_logic_vector(to_signed(1407,16));
        tmp(2021) := std_logic_vector(to_signed(1357,16));
        tmp(2022) := std_logic_vector(to_signed(1307,16));
        tmp(2023) := std_logic_vector(to_signed(1256,16));
        tmp(2024) := std_logic_vector(to_signed(1206,16));
        tmp(2025) := std_logic_vector(to_signed(1156,16));
        tmp(2026) := std_logic_vector(to_signed(1106,16));
        tmp(2027) := std_logic_vector(to_signed(1055,16));
        tmp(2028) := std_logic_vector(to_signed(1005,16));
        tmp(2029) := std_logic_vector(to_signed(955,16));
        tmp(2030) := std_logic_vector(to_signed(905,16));
        tmp(2031) := std_logic_vector(to_signed(854,16));
        tmp(2032) := std_logic_vector(to_signed(804,16));
        tmp(2033) := std_logic_vector(to_signed(754,16));
        tmp(2034) := std_logic_vector(to_signed(704,16));
        tmp(2035) := std_logic_vector(to_signed(653,16));
        tmp(2036) := std_logic_vector(to_signed(603,16));
        tmp(2037) := std_logic_vector(to_signed(553,16));
        tmp(2038) := std_logic_vector(to_signed(503,16));
        tmp(2039) := std_logic_vector(to_signed(452,16));
        tmp(2040) := std_logic_vector(to_signed(402,16));
        tmp(2041) := std_logic_vector(to_signed(352,16));
        tmp(2042) := std_logic_vector(to_signed(302,16));
        tmp(2043) := std_logic_vector(to_signed(251,16));
        tmp(2044) := std_logic_vector(to_signed(201,16));
        tmp(2045) := std_logic_vector(to_signed(151,16));
        tmp(2046) := std_logic_vector(to_signed(101,16));
        tmp(2047) := std_logic_vector(to_signed(50,16));
        tmp(2048) := std_logic_vector(to_signed(0,16));
        tmp(2049) := std_logic_vector(to_signed(-50,16));
        tmp(2050) := std_logic_vector(to_signed(-101,16));
        tmp(2051) := std_logic_vector(to_signed(-151,16));
        tmp(2052) := std_logic_vector(to_signed(-201,16));
        tmp(2053) := std_logic_vector(to_signed(-251,16));
        tmp(2054) := std_logic_vector(to_signed(-302,16));
        tmp(2055) := std_logic_vector(to_signed(-352,16));
        tmp(2056) := std_logic_vector(to_signed(-402,16));
        tmp(2057) := std_logic_vector(to_signed(-452,16));
        tmp(2058) := std_logic_vector(to_signed(-503,16));
        tmp(2059) := std_logic_vector(to_signed(-553,16));
        tmp(2060) := std_logic_vector(to_signed(-603,16));
        tmp(2061) := std_logic_vector(to_signed(-653,16));
        tmp(2062) := std_logic_vector(to_signed(-704,16));
        tmp(2063) := std_logic_vector(to_signed(-754,16));
        tmp(2064) := std_logic_vector(to_signed(-804,16));
        tmp(2065) := std_logic_vector(to_signed(-854,16));
        tmp(2066) := std_logic_vector(to_signed(-905,16));
        tmp(2067) := std_logic_vector(to_signed(-955,16));
        tmp(2068) := std_logic_vector(to_signed(-1005,16));
        tmp(2069) := std_logic_vector(to_signed(-1055,16));
        tmp(2070) := std_logic_vector(to_signed(-1106,16));
        tmp(2071) := std_logic_vector(to_signed(-1156,16));
        tmp(2072) := std_logic_vector(to_signed(-1206,16));
        tmp(2073) := std_logic_vector(to_signed(-1256,16));
        tmp(2074) := std_logic_vector(to_signed(-1307,16));
        tmp(2075) := std_logic_vector(to_signed(-1357,16));
        tmp(2076) := std_logic_vector(to_signed(-1407,16));
        tmp(2077) := std_logic_vector(to_signed(-1457,16));
        tmp(2078) := std_logic_vector(to_signed(-1507,16));
        tmp(2079) := std_logic_vector(to_signed(-1558,16));
        tmp(2080) := std_logic_vector(to_signed(-1608,16));
        tmp(2081) := std_logic_vector(to_signed(-1658,16));
        tmp(2082) := std_logic_vector(to_signed(-1708,16));
        tmp(2083) := std_logic_vector(to_signed(-1758,16));
        tmp(2084) := std_logic_vector(to_signed(-1809,16));
        tmp(2085) := std_logic_vector(to_signed(-1859,16));
        tmp(2086) := std_logic_vector(to_signed(-1909,16));
        tmp(2087) := std_logic_vector(to_signed(-1959,16));
        tmp(2088) := std_logic_vector(to_signed(-2009,16));
        tmp(2089) := std_logic_vector(to_signed(-2059,16));
        tmp(2090) := std_logic_vector(to_signed(-2110,16));
        tmp(2091) := std_logic_vector(to_signed(-2160,16));
        tmp(2092) := std_logic_vector(to_signed(-2210,16));
        tmp(2093) := std_logic_vector(to_signed(-2260,16));
        tmp(2094) := std_logic_vector(to_signed(-2310,16));
        tmp(2095) := std_logic_vector(to_signed(-2360,16));
        tmp(2096) := std_logic_vector(to_signed(-2410,16));
        tmp(2097) := std_logic_vector(to_signed(-2461,16));
        tmp(2098) := std_logic_vector(to_signed(-2511,16));
        tmp(2099) := std_logic_vector(to_signed(-2561,16));
        tmp(2100) := std_logic_vector(to_signed(-2611,16));
        tmp(2101) := std_logic_vector(to_signed(-2661,16));
        tmp(2102) := std_logic_vector(to_signed(-2711,16));
        tmp(2103) := std_logic_vector(to_signed(-2761,16));
        tmp(2104) := std_logic_vector(to_signed(-2811,16));
        tmp(2105) := std_logic_vector(to_signed(-2861,16));
        tmp(2106) := std_logic_vector(to_signed(-2911,16));
        tmp(2107) := std_logic_vector(to_signed(-2962,16));
        tmp(2108) := std_logic_vector(to_signed(-3012,16));
        tmp(2109) := std_logic_vector(to_signed(-3062,16));
        tmp(2110) := std_logic_vector(to_signed(-3112,16));
        tmp(2111) := std_logic_vector(to_signed(-3162,16));
        tmp(2112) := std_logic_vector(to_signed(-3212,16));
        tmp(2113) := std_logic_vector(to_signed(-3262,16));
        tmp(2114) := std_logic_vector(to_signed(-3312,16));
        tmp(2115) := std_logic_vector(to_signed(-3362,16));
        tmp(2116) := std_logic_vector(to_signed(-3412,16));
        tmp(2117) := std_logic_vector(to_signed(-3462,16));
        tmp(2118) := std_logic_vector(to_signed(-3512,16));
        tmp(2119) := std_logic_vector(to_signed(-3562,16));
        tmp(2120) := std_logic_vector(to_signed(-3612,16));
        tmp(2121) := std_logic_vector(to_signed(-3662,16));
        tmp(2122) := std_logic_vector(to_signed(-3712,16));
        tmp(2123) := std_logic_vector(to_signed(-3761,16));
        tmp(2124) := std_logic_vector(to_signed(-3811,16));
        tmp(2125) := std_logic_vector(to_signed(-3861,16));
        tmp(2126) := std_logic_vector(to_signed(-3911,16));
        tmp(2127) := std_logic_vector(to_signed(-3961,16));
        tmp(2128) := std_logic_vector(to_signed(-4011,16));
        tmp(2129) := std_logic_vector(to_signed(-4061,16));
        tmp(2130) := std_logic_vector(to_signed(-4111,16));
        tmp(2131) := std_logic_vector(to_signed(-4161,16));
        tmp(2132) := std_logic_vector(to_signed(-4210,16));
        tmp(2133) := std_logic_vector(to_signed(-4260,16));
        tmp(2134) := std_logic_vector(to_signed(-4310,16));
        tmp(2135) := std_logic_vector(to_signed(-4360,16));
        tmp(2136) := std_logic_vector(to_signed(-4410,16));
        tmp(2137) := std_logic_vector(to_signed(-4460,16));
        tmp(2138) := std_logic_vector(to_signed(-4509,16));
        tmp(2139) := std_logic_vector(to_signed(-4559,16));
        tmp(2140) := std_logic_vector(to_signed(-4609,16));
        tmp(2141) := std_logic_vector(to_signed(-4659,16));
        tmp(2142) := std_logic_vector(to_signed(-4708,16));
        tmp(2143) := std_logic_vector(to_signed(-4758,16));
        tmp(2144) := std_logic_vector(to_signed(-4808,16));
        tmp(2145) := std_logic_vector(to_signed(-4858,16));
        tmp(2146) := std_logic_vector(to_signed(-4907,16));
        tmp(2147) := std_logic_vector(to_signed(-4957,16));
        tmp(2148) := std_logic_vector(to_signed(-5007,16));
        tmp(2149) := std_logic_vector(to_signed(-5056,16));
        tmp(2150) := std_logic_vector(to_signed(-5106,16));
        tmp(2151) := std_logic_vector(to_signed(-5156,16));
        tmp(2152) := std_logic_vector(to_signed(-5205,16));
        tmp(2153) := std_logic_vector(to_signed(-5255,16));
        tmp(2154) := std_logic_vector(to_signed(-5305,16));
        tmp(2155) := std_logic_vector(to_signed(-5354,16));
        tmp(2156) := std_logic_vector(to_signed(-5404,16));
        tmp(2157) := std_logic_vector(to_signed(-5453,16));
        tmp(2158) := std_logic_vector(to_signed(-5503,16));
        tmp(2159) := std_logic_vector(to_signed(-5552,16));
        tmp(2160) := std_logic_vector(to_signed(-5602,16));
        tmp(2161) := std_logic_vector(to_signed(-5651,16));
        tmp(2162) := std_logic_vector(to_signed(-5701,16));
        tmp(2163) := std_logic_vector(to_signed(-5750,16));
        tmp(2164) := std_logic_vector(to_signed(-5800,16));
        tmp(2165) := std_logic_vector(to_signed(-5849,16));
        tmp(2166) := std_logic_vector(to_signed(-5899,16));
        tmp(2167) := std_logic_vector(to_signed(-5948,16));
        tmp(2168) := std_logic_vector(to_signed(-5998,16));
        tmp(2169) := std_logic_vector(to_signed(-6047,16));
        tmp(2170) := std_logic_vector(to_signed(-6096,16));
        tmp(2171) := std_logic_vector(to_signed(-6146,16));
        tmp(2172) := std_logic_vector(to_signed(-6195,16));
        tmp(2173) := std_logic_vector(to_signed(-6245,16));
        tmp(2174) := std_logic_vector(to_signed(-6294,16));
        tmp(2175) := std_logic_vector(to_signed(-6343,16));
        tmp(2176) := std_logic_vector(to_signed(-6393,16));
        tmp(2177) := std_logic_vector(to_signed(-6442,16));
        tmp(2178) := std_logic_vector(to_signed(-6491,16));
        tmp(2179) := std_logic_vector(to_signed(-6540,16));
        tmp(2180) := std_logic_vector(to_signed(-6590,16));
        tmp(2181) := std_logic_vector(to_signed(-6639,16));
        tmp(2182) := std_logic_vector(to_signed(-6688,16));
        tmp(2183) := std_logic_vector(to_signed(-6737,16));
        tmp(2184) := std_logic_vector(to_signed(-6786,16));
        tmp(2185) := std_logic_vector(to_signed(-6836,16));
        tmp(2186) := std_logic_vector(to_signed(-6885,16));
        tmp(2187) := std_logic_vector(to_signed(-6934,16));
        tmp(2188) := std_logic_vector(to_signed(-6983,16));
        tmp(2189) := std_logic_vector(to_signed(-7032,16));
        tmp(2190) := std_logic_vector(to_signed(-7081,16));
        tmp(2191) := std_logic_vector(to_signed(-7130,16));
        tmp(2192) := std_logic_vector(to_signed(-7179,16));
        tmp(2193) := std_logic_vector(to_signed(-7228,16));
        tmp(2194) := std_logic_vector(to_signed(-7277,16));
        tmp(2195) := std_logic_vector(to_signed(-7326,16));
        tmp(2196) := std_logic_vector(to_signed(-7375,16));
        tmp(2197) := std_logic_vector(to_signed(-7424,16));
        tmp(2198) := std_logic_vector(to_signed(-7473,16));
        tmp(2199) := std_logic_vector(to_signed(-7522,16));
        tmp(2200) := std_logic_vector(to_signed(-7571,16));
        tmp(2201) := std_logic_vector(to_signed(-7620,16));
        tmp(2202) := std_logic_vector(to_signed(-7669,16));
        tmp(2203) := std_logic_vector(to_signed(-7718,16));
        tmp(2204) := std_logic_vector(to_signed(-7767,16));
        tmp(2205) := std_logic_vector(to_signed(-7815,16));
        tmp(2206) := std_logic_vector(to_signed(-7864,16));
        tmp(2207) := std_logic_vector(to_signed(-7913,16));
        tmp(2208) := std_logic_vector(to_signed(-7962,16));
        tmp(2209) := std_logic_vector(to_signed(-8010,16));
        tmp(2210) := std_logic_vector(to_signed(-8059,16));
        tmp(2211) := std_logic_vector(to_signed(-8108,16));
        tmp(2212) := std_logic_vector(to_signed(-8157,16));
        tmp(2213) := std_logic_vector(to_signed(-8205,16));
        tmp(2214) := std_logic_vector(to_signed(-8254,16));
        tmp(2215) := std_logic_vector(to_signed(-8303,16));
        tmp(2216) := std_logic_vector(to_signed(-8351,16));
        tmp(2217) := std_logic_vector(to_signed(-8400,16));
        tmp(2218) := std_logic_vector(to_signed(-8448,16));
        tmp(2219) := std_logic_vector(to_signed(-8497,16));
        tmp(2220) := std_logic_vector(to_signed(-8545,16));
        tmp(2221) := std_logic_vector(to_signed(-8594,16));
        tmp(2222) := std_logic_vector(to_signed(-8642,16));
        tmp(2223) := std_logic_vector(to_signed(-8691,16));
        tmp(2224) := std_logic_vector(to_signed(-8739,16));
        tmp(2225) := std_logic_vector(to_signed(-8788,16));
        tmp(2226) := std_logic_vector(to_signed(-8836,16));
        tmp(2227) := std_logic_vector(to_signed(-8885,16));
        tmp(2228) := std_logic_vector(to_signed(-8933,16));
        tmp(2229) := std_logic_vector(to_signed(-8981,16));
        tmp(2230) := std_logic_vector(to_signed(-9030,16));
        tmp(2231) := std_logic_vector(to_signed(-9078,16));
        tmp(2232) := std_logic_vector(to_signed(-9126,16));
        tmp(2233) := std_logic_vector(to_signed(-9175,16));
        tmp(2234) := std_logic_vector(to_signed(-9223,16));
        tmp(2235) := std_logic_vector(to_signed(-9271,16));
        tmp(2236) := std_logic_vector(to_signed(-9319,16));
        tmp(2237) := std_logic_vector(to_signed(-9367,16));
        tmp(2238) := std_logic_vector(to_signed(-9416,16));
        tmp(2239) := std_logic_vector(to_signed(-9464,16));
        tmp(2240) := std_logic_vector(to_signed(-9512,16));
        tmp(2241) := std_logic_vector(to_signed(-9560,16));
        tmp(2242) := std_logic_vector(to_signed(-9608,16));
        tmp(2243) := std_logic_vector(to_signed(-9656,16));
        tmp(2244) := std_logic_vector(to_signed(-9704,16));
        tmp(2245) := std_logic_vector(to_signed(-9752,16));
        tmp(2246) := std_logic_vector(to_signed(-9800,16));
        tmp(2247) := std_logic_vector(to_signed(-9848,16));
        tmp(2248) := std_logic_vector(to_signed(-9896,16));
        tmp(2249) := std_logic_vector(to_signed(-9944,16));
        tmp(2250) := std_logic_vector(to_signed(-9992,16));
        tmp(2251) := std_logic_vector(to_signed(-10039,16));
        tmp(2252) := std_logic_vector(to_signed(-10087,16));
        tmp(2253) := std_logic_vector(to_signed(-10135,16));
        tmp(2254) := std_logic_vector(to_signed(-10183,16));
        tmp(2255) := std_logic_vector(to_signed(-10231,16));
        tmp(2256) := std_logic_vector(to_signed(-10278,16));
        tmp(2257) := std_logic_vector(to_signed(-10326,16));
        tmp(2258) := std_logic_vector(to_signed(-10374,16));
        tmp(2259) := std_logic_vector(to_signed(-10421,16));
        tmp(2260) := std_logic_vector(to_signed(-10469,16));
        tmp(2261) := std_logic_vector(to_signed(-10517,16));
        tmp(2262) := std_logic_vector(to_signed(-10564,16));
        tmp(2263) := std_logic_vector(to_signed(-10612,16));
        tmp(2264) := std_logic_vector(to_signed(-10659,16));
        tmp(2265) := std_logic_vector(to_signed(-10707,16));
        tmp(2266) := std_logic_vector(to_signed(-10754,16));
        tmp(2267) := std_logic_vector(to_signed(-10802,16));
        tmp(2268) := std_logic_vector(to_signed(-10849,16));
        tmp(2269) := std_logic_vector(to_signed(-10897,16));
        tmp(2270) := std_logic_vector(to_signed(-10944,16));
        tmp(2271) := std_logic_vector(to_signed(-10992,16));
        tmp(2272) := std_logic_vector(to_signed(-11039,16));
        tmp(2273) := std_logic_vector(to_signed(-11086,16));
        tmp(2274) := std_logic_vector(to_signed(-11133,16));
        tmp(2275) := std_logic_vector(to_signed(-11181,16));
        tmp(2276) := std_logic_vector(to_signed(-11228,16));
        tmp(2277) := std_logic_vector(to_signed(-11275,16));
        tmp(2278) := std_logic_vector(to_signed(-11322,16));
        tmp(2279) := std_logic_vector(to_signed(-11370,16));
        tmp(2280) := std_logic_vector(to_signed(-11417,16));
        tmp(2281) := std_logic_vector(to_signed(-11464,16));
        tmp(2282) := std_logic_vector(to_signed(-11511,16));
        tmp(2283) := std_logic_vector(to_signed(-11558,16));
        tmp(2284) := std_logic_vector(to_signed(-11605,16));
        tmp(2285) := std_logic_vector(to_signed(-11652,16));
        tmp(2286) := std_logic_vector(to_signed(-11699,16));
        tmp(2287) := std_logic_vector(to_signed(-11746,16));
        tmp(2288) := std_logic_vector(to_signed(-11793,16));
        tmp(2289) := std_logic_vector(to_signed(-11840,16));
        tmp(2290) := std_logic_vector(to_signed(-11886,16));
        tmp(2291) := std_logic_vector(to_signed(-11933,16));
        tmp(2292) := std_logic_vector(to_signed(-11980,16));
        tmp(2293) := std_logic_vector(to_signed(-12027,16));
        tmp(2294) := std_logic_vector(to_signed(-12074,16));
        tmp(2295) := std_logic_vector(to_signed(-12120,16));
        tmp(2296) := std_logic_vector(to_signed(-12167,16));
        tmp(2297) := std_logic_vector(to_signed(-12214,16));
        tmp(2298) := std_logic_vector(to_signed(-12260,16));
        tmp(2299) := std_logic_vector(to_signed(-12307,16));
        tmp(2300) := std_logic_vector(to_signed(-12353,16));
        tmp(2301) := std_logic_vector(to_signed(-12400,16));
        tmp(2302) := std_logic_vector(to_signed(-12446,16));
        tmp(2303) := std_logic_vector(to_signed(-12493,16));
        tmp(2304) := std_logic_vector(to_signed(-12539,16));
        tmp(2305) := std_logic_vector(to_signed(-12586,16));
        tmp(2306) := std_logic_vector(to_signed(-12632,16));
        tmp(2307) := std_logic_vector(to_signed(-12679,16));
        tmp(2308) := std_logic_vector(to_signed(-12725,16));
        tmp(2309) := std_logic_vector(to_signed(-12771,16));
        tmp(2310) := std_logic_vector(to_signed(-12817,16));
        tmp(2311) := std_logic_vector(to_signed(-12864,16));
        tmp(2312) := std_logic_vector(to_signed(-12910,16));
        tmp(2313) := std_logic_vector(to_signed(-12956,16));
        tmp(2314) := std_logic_vector(to_signed(-13002,16));
        tmp(2315) := std_logic_vector(to_signed(-13048,16));
        tmp(2316) := std_logic_vector(to_signed(-13094,16));
        tmp(2317) := std_logic_vector(to_signed(-13141,16));
        tmp(2318) := std_logic_vector(to_signed(-13187,16));
        tmp(2319) := std_logic_vector(to_signed(-13233,16));
        tmp(2320) := std_logic_vector(to_signed(-13279,16));
        tmp(2321) := std_logic_vector(to_signed(-13324,16));
        tmp(2322) := std_logic_vector(to_signed(-13370,16));
        tmp(2323) := std_logic_vector(to_signed(-13416,16));
        tmp(2324) := std_logic_vector(to_signed(-13462,16));
        tmp(2325) := std_logic_vector(to_signed(-13508,16));
        tmp(2326) := std_logic_vector(to_signed(-13554,16));
        tmp(2327) := std_logic_vector(to_signed(-13599,16));
        tmp(2328) := std_logic_vector(to_signed(-13645,16));
        tmp(2329) := std_logic_vector(to_signed(-13691,16));
        tmp(2330) := std_logic_vector(to_signed(-13736,16));
        tmp(2331) := std_logic_vector(to_signed(-13782,16));
        tmp(2332) := std_logic_vector(to_signed(-13828,16));
        tmp(2333) := std_logic_vector(to_signed(-13873,16));
        tmp(2334) := std_logic_vector(to_signed(-13919,16));
        tmp(2335) := std_logic_vector(to_signed(-13964,16));
        tmp(2336) := std_logic_vector(to_signed(-14010,16));
        tmp(2337) := std_logic_vector(to_signed(-14055,16));
        tmp(2338) := std_logic_vector(to_signed(-14101,16));
        tmp(2339) := std_logic_vector(to_signed(-14146,16));
        tmp(2340) := std_logic_vector(to_signed(-14191,16));
        tmp(2341) := std_logic_vector(to_signed(-14236,16));
        tmp(2342) := std_logic_vector(to_signed(-14282,16));
        tmp(2343) := std_logic_vector(to_signed(-14327,16));
        tmp(2344) := std_logic_vector(to_signed(-14372,16));
        tmp(2345) := std_logic_vector(to_signed(-14417,16));
        tmp(2346) := std_logic_vector(to_signed(-14462,16));
        tmp(2347) := std_logic_vector(to_signed(-14507,16));
        tmp(2348) := std_logic_vector(to_signed(-14553,16));
        tmp(2349) := std_logic_vector(to_signed(-14598,16));
        tmp(2350) := std_logic_vector(to_signed(-14643,16));
        tmp(2351) := std_logic_vector(to_signed(-14688,16));
        tmp(2352) := std_logic_vector(to_signed(-14732,16));
        tmp(2353) := std_logic_vector(to_signed(-14777,16));
        tmp(2354) := std_logic_vector(to_signed(-14822,16));
        tmp(2355) := std_logic_vector(to_signed(-14867,16));
        tmp(2356) := std_logic_vector(to_signed(-14912,16));
        tmp(2357) := std_logic_vector(to_signed(-14956,16));
        tmp(2358) := std_logic_vector(to_signed(-15001,16));
        tmp(2359) := std_logic_vector(to_signed(-15046,16));
        tmp(2360) := std_logic_vector(to_signed(-15090,16));
        tmp(2361) := std_logic_vector(to_signed(-15135,16));
        tmp(2362) := std_logic_vector(to_signed(-15180,16));
        tmp(2363) := std_logic_vector(to_signed(-15224,16));
        tmp(2364) := std_logic_vector(to_signed(-15269,16));
        tmp(2365) := std_logic_vector(to_signed(-15313,16));
        tmp(2366) := std_logic_vector(to_signed(-15358,16));
        tmp(2367) := std_logic_vector(to_signed(-15402,16));
        tmp(2368) := std_logic_vector(to_signed(-15446,16));
        tmp(2369) := std_logic_vector(to_signed(-15491,16));
        tmp(2370) := std_logic_vector(to_signed(-15535,16));
        tmp(2371) := std_logic_vector(to_signed(-15579,16));
        tmp(2372) := std_logic_vector(to_signed(-15623,16));
        tmp(2373) := std_logic_vector(to_signed(-15667,16));
        tmp(2374) := std_logic_vector(to_signed(-15712,16));
        tmp(2375) := std_logic_vector(to_signed(-15756,16));
        tmp(2376) := std_logic_vector(to_signed(-15800,16));
        tmp(2377) := std_logic_vector(to_signed(-15844,16));
        tmp(2378) := std_logic_vector(to_signed(-15888,16));
        tmp(2379) := std_logic_vector(to_signed(-15932,16));
        tmp(2380) := std_logic_vector(to_signed(-15976,16));
        tmp(2381) := std_logic_vector(to_signed(-16019,16));
        tmp(2382) := std_logic_vector(to_signed(-16063,16));
        tmp(2383) := std_logic_vector(to_signed(-16107,16));
        tmp(2384) := std_logic_vector(to_signed(-16151,16));
        tmp(2385) := std_logic_vector(to_signed(-16195,16));
        tmp(2386) := std_logic_vector(to_signed(-16238,16));
        tmp(2387) := std_logic_vector(to_signed(-16282,16));
        tmp(2388) := std_logic_vector(to_signed(-16325,16));
        tmp(2389) := std_logic_vector(to_signed(-16369,16));
        tmp(2390) := std_logic_vector(to_signed(-16413,16));
        tmp(2391) := std_logic_vector(to_signed(-16456,16));
        tmp(2392) := std_logic_vector(to_signed(-16499,16));
        tmp(2393) := std_logic_vector(to_signed(-16543,16));
        tmp(2394) := std_logic_vector(to_signed(-16586,16));
        tmp(2395) := std_logic_vector(to_signed(-16630,16));
        tmp(2396) := std_logic_vector(to_signed(-16673,16));
        tmp(2397) := std_logic_vector(to_signed(-16716,16));
        tmp(2398) := std_logic_vector(to_signed(-16759,16));
        tmp(2399) := std_logic_vector(to_signed(-16802,16));
        tmp(2400) := std_logic_vector(to_signed(-16846,16));
        tmp(2401) := std_logic_vector(to_signed(-16889,16));
        tmp(2402) := std_logic_vector(to_signed(-16932,16));
        tmp(2403) := std_logic_vector(to_signed(-16975,16));
        tmp(2404) := std_logic_vector(to_signed(-17018,16));
        tmp(2405) := std_logic_vector(to_signed(-17061,16));
        tmp(2406) := std_logic_vector(to_signed(-17104,16));
        tmp(2407) := std_logic_vector(to_signed(-17146,16));
        tmp(2408) := std_logic_vector(to_signed(-17189,16));
        tmp(2409) := std_logic_vector(to_signed(-17232,16));
        tmp(2410) := std_logic_vector(to_signed(-17275,16));
        tmp(2411) := std_logic_vector(to_signed(-17317,16));
        tmp(2412) := std_logic_vector(to_signed(-17360,16));
        tmp(2413) := std_logic_vector(to_signed(-17403,16));
        tmp(2414) := std_logic_vector(to_signed(-17445,16));
        tmp(2415) := std_logic_vector(to_signed(-17488,16));
        tmp(2416) := std_logic_vector(to_signed(-17530,16));
        tmp(2417) := std_logic_vector(to_signed(-17573,16));
        tmp(2418) := std_logic_vector(to_signed(-17615,16));
        tmp(2419) := std_logic_vector(to_signed(-17657,16));
        tmp(2420) := std_logic_vector(to_signed(-17700,16));
        tmp(2421) := std_logic_vector(to_signed(-17742,16));
        tmp(2422) := std_logic_vector(to_signed(-17784,16));
        tmp(2423) := std_logic_vector(to_signed(-17827,16));
        tmp(2424) := std_logic_vector(to_signed(-17869,16));
        tmp(2425) := std_logic_vector(to_signed(-17911,16));
        tmp(2426) := std_logic_vector(to_signed(-17953,16));
        tmp(2427) := std_logic_vector(to_signed(-17995,16));
        tmp(2428) := std_logic_vector(to_signed(-18037,16));
        tmp(2429) := std_logic_vector(to_signed(-18079,16));
        tmp(2430) := std_logic_vector(to_signed(-18121,16));
        tmp(2431) := std_logic_vector(to_signed(-18163,16));
        tmp(2432) := std_logic_vector(to_signed(-18204,16));
        tmp(2433) := std_logic_vector(to_signed(-18246,16));
        tmp(2434) := std_logic_vector(to_signed(-18288,16));
        tmp(2435) := std_logic_vector(to_signed(-18330,16));
        tmp(2436) := std_logic_vector(to_signed(-18371,16));
        tmp(2437) := std_logic_vector(to_signed(-18413,16));
        tmp(2438) := std_logic_vector(to_signed(-18454,16));
        tmp(2439) := std_logic_vector(to_signed(-18496,16));
        tmp(2440) := std_logic_vector(to_signed(-18537,16));
        tmp(2441) := std_logic_vector(to_signed(-18579,16));
        tmp(2442) := std_logic_vector(to_signed(-18620,16));
        tmp(2443) := std_logic_vector(to_signed(-18661,16));
        tmp(2444) := std_logic_vector(to_signed(-18703,16));
        tmp(2445) := std_logic_vector(to_signed(-18744,16));
        tmp(2446) := std_logic_vector(to_signed(-18785,16));
        tmp(2447) := std_logic_vector(to_signed(-18826,16));
        tmp(2448) := std_logic_vector(to_signed(-18868,16));
        tmp(2449) := std_logic_vector(to_signed(-18909,16));
        tmp(2450) := std_logic_vector(to_signed(-18950,16));
        tmp(2451) := std_logic_vector(to_signed(-18991,16));
        tmp(2452) := std_logic_vector(to_signed(-19032,16));
        tmp(2453) := std_logic_vector(to_signed(-19072,16));
        tmp(2454) := std_logic_vector(to_signed(-19113,16));
        tmp(2455) := std_logic_vector(to_signed(-19154,16));
        tmp(2456) := std_logic_vector(to_signed(-19195,16));
        tmp(2457) := std_logic_vector(to_signed(-19236,16));
        tmp(2458) := std_logic_vector(to_signed(-19276,16));
        tmp(2459) := std_logic_vector(to_signed(-19317,16));
        tmp(2460) := std_logic_vector(to_signed(-19357,16));
        tmp(2461) := std_logic_vector(to_signed(-19398,16));
        tmp(2462) := std_logic_vector(to_signed(-19438,16));
        tmp(2463) := std_logic_vector(to_signed(-19479,16));
        tmp(2464) := std_logic_vector(to_signed(-19519,16));
        tmp(2465) := std_logic_vector(to_signed(-19560,16));
        tmp(2466) := std_logic_vector(to_signed(-19600,16));
        tmp(2467) := std_logic_vector(to_signed(-19640,16));
        tmp(2468) := std_logic_vector(to_signed(-19680,16));
        tmp(2469) := std_logic_vector(to_signed(-19721,16));
        tmp(2470) := std_logic_vector(to_signed(-19761,16));
        tmp(2471) := std_logic_vector(to_signed(-19801,16));
        tmp(2472) := std_logic_vector(to_signed(-19841,16));
        tmp(2473) := std_logic_vector(to_signed(-19881,16));
        tmp(2474) := std_logic_vector(to_signed(-19921,16));
        tmp(2475) := std_logic_vector(to_signed(-19961,16));
        tmp(2476) := std_logic_vector(to_signed(-20000,16));
        tmp(2477) := std_logic_vector(to_signed(-20040,16));
        tmp(2478) := std_logic_vector(to_signed(-20080,16));
        tmp(2479) := std_logic_vector(to_signed(-20120,16));
        tmp(2480) := std_logic_vector(to_signed(-20159,16));
        tmp(2481) := std_logic_vector(to_signed(-20199,16));
        tmp(2482) := std_logic_vector(to_signed(-20238,16));
        tmp(2483) := std_logic_vector(to_signed(-20278,16));
        tmp(2484) := std_logic_vector(to_signed(-20317,16));
        tmp(2485) := std_logic_vector(to_signed(-20357,16));
        tmp(2486) := std_logic_vector(to_signed(-20396,16));
        tmp(2487) := std_logic_vector(to_signed(-20436,16));
        tmp(2488) := std_logic_vector(to_signed(-20475,16));
        tmp(2489) := std_logic_vector(to_signed(-20514,16));
        tmp(2490) := std_logic_vector(to_signed(-20553,16));
        tmp(2491) := std_logic_vector(to_signed(-20592,16));
        tmp(2492) := std_logic_vector(to_signed(-20631,16));
        tmp(2493) := std_logic_vector(to_signed(-20670,16));
        tmp(2494) := std_logic_vector(to_signed(-20709,16));
        tmp(2495) := std_logic_vector(to_signed(-20748,16));
        tmp(2496) := std_logic_vector(to_signed(-20787,16));
        tmp(2497) := std_logic_vector(to_signed(-20826,16));
        tmp(2498) := std_logic_vector(to_signed(-20865,16));
        tmp(2499) := std_logic_vector(to_signed(-20904,16));
        tmp(2500) := std_logic_vector(to_signed(-20942,16));
        tmp(2501) := std_logic_vector(to_signed(-20981,16));
        tmp(2502) := std_logic_vector(to_signed(-21019,16));
        tmp(2503) := std_logic_vector(to_signed(-21058,16));
        tmp(2504) := std_logic_vector(to_signed(-21096,16));
        tmp(2505) := std_logic_vector(to_signed(-21135,16));
        tmp(2506) := std_logic_vector(to_signed(-21173,16));
        tmp(2507) := std_logic_vector(to_signed(-21212,16));
        tmp(2508) := std_logic_vector(to_signed(-21250,16));
        tmp(2509) := std_logic_vector(to_signed(-21288,16));
        tmp(2510) := std_logic_vector(to_signed(-21326,16));
        tmp(2511) := std_logic_vector(to_signed(-21364,16));
        tmp(2512) := std_logic_vector(to_signed(-21403,16));
        tmp(2513) := std_logic_vector(to_signed(-21441,16));
        tmp(2514) := std_logic_vector(to_signed(-21479,16));
        tmp(2515) := std_logic_vector(to_signed(-21516,16));
        tmp(2516) := std_logic_vector(to_signed(-21554,16));
        tmp(2517) := std_logic_vector(to_signed(-21592,16));
        tmp(2518) := std_logic_vector(to_signed(-21630,16));
        tmp(2519) := std_logic_vector(to_signed(-21668,16));
        tmp(2520) := std_logic_vector(to_signed(-21705,16));
        tmp(2521) := std_logic_vector(to_signed(-21743,16));
        tmp(2522) := std_logic_vector(to_signed(-21781,16));
        tmp(2523) := std_logic_vector(to_signed(-21818,16));
        tmp(2524) := std_logic_vector(to_signed(-21856,16));
        tmp(2525) := std_logic_vector(to_signed(-21893,16));
        tmp(2526) := std_logic_vector(to_signed(-21930,16));
        tmp(2527) := std_logic_vector(to_signed(-21968,16));
        tmp(2528) := std_logic_vector(to_signed(-22005,16));
        tmp(2529) := std_logic_vector(to_signed(-22042,16));
        tmp(2530) := std_logic_vector(to_signed(-22079,16));
        tmp(2531) := std_logic_vector(to_signed(-22116,16));
        tmp(2532) := std_logic_vector(to_signed(-22154,16));
        tmp(2533) := std_logic_vector(to_signed(-22191,16));
        tmp(2534) := std_logic_vector(to_signed(-22227,16));
        tmp(2535) := std_logic_vector(to_signed(-22264,16));
        tmp(2536) := std_logic_vector(to_signed(-22301,16));
        tmp(2537) := std_logic_vector(to_signed(-22338,16));
        tmp(2538) := std_logic_vector(to_signed(-22375,16));
        tmp(2539) := std_logic_vector(to_signed(-22411,16));
        tmp(2540) := std_logic_vector(to_signed(-22448,16));
        tmp(2541) := std_logic_vector(to_signed(-22485,16));
        tmp(2542) := std_logic_vector(to_signed(-22521,16));
        tmp(2543) := std_logic_vector(to_signed(-22558,16));
        tmp(2544) := std_logic_vector(to_signed(-22594,16));
        tmp(2545) := std_logic_vector(to_signed(-22631,16));
        tmp(2546) := std_logic_vector(to_signed(-22667,16));
        tmp(2547) := std_logic_vector(to_signed(-22703,16));
        tmp(2548) := std_logic_vector(to_signed(-22739,16));
        tmp(2549) := std_logic_vector(to_signed(-22776,16));
        tmp(2550) := std_logic_vector(to_signed(-22812,16));
        tmp(2551) := std_logic_vector(to_signed(-22848,16));
        tmp(2552) := std_logic_vector(to_signed(-22884,16));
        tmp(2553) := std_logic_vector(to_signed(-22920,16));
        tmp(2554) := std_logic_vector(to_signed(-22956,16));
        tmp(2555) := std_logic_vector(to_signed(-22991,16));
        tmp(2556) := std_logic_vector(to_signed(-23027,16));
        tmp(2557) := std_logic_vector(to_signed(-23063,16));
        tmp(2558) := std_logic_vector(to_signed(-23099,16));
        tmp(2559) := std_logic_vector(to_signed(-23134,16));
        tmp(2560) := std_logic_vector(to_signed(-23170,16));
        tmp(2561) := std_logic_vector(to_signed(-23205,16));
        tmp(2562) := std_logic_vector(to_signed(-23241,16));
        tmp(2563) := std_logic_vector(to_signed(-23276,16));
        tmp(2564) := std_logic_vector(to_signed(-23311,16));
        tmp(2565) := std_logic_vector(to_signed(-23347,16));
        tmp(2566) := std_logic_vector(to_signed(-23382,16));
        tmp(2567) := std_logic_vector(to_signed(-23417,16));
        tmp(2568) := std_logic_vector(to_signed(-23452,16));
        tmp(2569) := std_logic_vector(to_signed(-23487,16));
        tmp(2570) := std_logic_vector(to_signed(-23522,16));
        tmp(2571) := std_logic_vector(to_signed(-23557,16));
        tmp(2572) := std_logic_vector(to_signed(-23592,16));
        tmp(2573) := std_logic_vector(to_signed(-23627,16));
        tmp(2574) := std_logic_vector(to_signed(-23662,16));
        tmp(2575) := std_logic_vector(to_signed(-23697,16));
        tmp(2576) := std_logic_vector(to_signed(-23731,16));
        tmp(2577) := std_logic_vector(to_signed(-23766,16));
        tmp(2578) := std_logic_vector(to_signed(-23801,16));
        tmp(2579) := std_logic_vector(to_signed(-23835,16));
        tmp(2580) := std_logic_vector(to_signed(-23870,16));
        tmp(2581) := std_logic_vector(to_signed(-23904,16));
        tmp(2582) := std_logic_vector(to_signed(-23938,16));
        tmp(2583) := std_logic_vector(to_signed(-23973,16));
        tmp(2584) := std_logic_vector(to_signed(-24007,16));
        tmp(2585) := std_logic_vector(to_signed(-24041,16));
        tmp(2586) := std_logic_vector(to_signed(-24075,16));
        tmp(2587) := std_logic_vector(to_signed(-24109,16));
        tmp(2588) := std_logic_vector(to_signed(-24143,16));
        tmp(2589) := std_logic_vector(to_signed(-24177,16));
        tmp(2590) := std_logic_vector(to_signed(-24211,16));
        tmp(2591) := std_logic_vector(to_signed(-24245,16));
        tmp(2592) := std_logic_vector(to_signed(-24279,16));
        tmp(2593) := std_logic_vector(to_signed(-24312,16));
        tmp(2594) := std_logic_vector(to_signed(-24346,16));
        tmp(2595) := std_logic_vector(to_signed(-24380,16));
        tmp(2596) := std_logic_vector(to_signed(-24413,16));
        tmp(2597) := std_logic_vector(to_signed(-24447,16));
        tmp(2598) := std_logic_vector(to_signed(-24480,16));
        tmp(2599) := std_logic_vector(to_signed(-24514,16));
        tmp(2600) := std_logic_vector(to_signed(-24547,16));
        tmp(2601) := std_logic_vector(to_signed(-24580,16));
        tmp(2602) := std_logic_vector(to_signed(-24613,16));
        tmp(2603) := std_logic_vector(to_signed(-24647,16));
        tmp(2604) := std_logic_vector(to_signed(-24680,16));
        tmp(2605) := std_logic_vector(to_signed(-24713,16));
        tmp(2606) := std_logic_vector(to_signed(-24746,16));
        tmp(2607) := std_logic_vector(to_signed(-24779,16));
        tmp(2608) := std_logic_vector(to_signed(-24811,16));
        tmp(2609) := std_logic_vector(to_signed(-24844,16));
        tmp(2610) := std_logic_vector(to_signed(-24877,16));
        tmp(2611) := std_logic_vector(to_signed(-24910,16));
        tmp(2612) := std_logic_vector(to_signed(-24942,16));
        tmp(2613) := std_logic_vector(to_signed(-24975,16));
        tmp(2614) := std_logic_vector(to_signed(-25007,16));
        tmp(2615) := std_logic_vector(to_signed(-25040,16));
        tmp(2616) := std_logic_vector(to_signed(-25072,16));
        tmp(2617) := std_logic_vector(to_signed(-25105,16));
        tmp(2618) := std_logic_vector(to_signed(-25137,16));
        tmp(2619) := std_logic_vector(to_signed(-25169,16));
        tmp(2620) := std_logic_vector(to_signed(-25201,16));
        tmp(2621) := std_logic_vector(to_signed(-25233,16));
        tmp(2622) := std_logic_vector(to_signed(-25265,16));
        tmp(2623) := std_logic_vector(to_signed(-25297,16));
        tmp(2624) := std_logic_vector(to_signed(-25329,16));
        tmp(2625) := std_logic_vector(to_signed(-25361,16));
        tmp(2626) := std_logic_vector(to_signed(-25393,16));
        tmp(2627) := std_logic_vector(to_signed(-25425,16));
        tmp(2628) := std_logic_vector(to_signed(-25456,16));
        tmp(2629) := std_logic_vector(to_signed(-25488,16));
        tmp(2630) := std_logic_vector(to_signed(-25519,16));
        tmp(2631) := std_logic_vector(to_signed(-25551,16));
        tmp(2632) := std_logic_vector(to_signed(-25582,16));
        tmp(2633) := std_logic_vector(to_signed(-25614,16));
        tmp(2634) := std_logic_vector(to_signed(-25645,16));
        tmp(2635) := std_logic_vector(to_signed(-25676,16));
        tmp(2636) := std_logic_vector(to_signed(-25708,16));
        tmp(2637) := std_logic_vector(to_signed(-25739,16));
        tmp(2638) := std_logic_vector(to_signed(-25770,16));
        tmp(2639) := std_logic_vector(to_signed(-25801,16));
        tmp(2640) := std_logic_vector(to_signed(-25832,16));
        tmp(2641) := std_logic_vector(to_signed(-25863,16));
        tmp(2642) := std_logic_vector(to_signed(-25893,16));
        tmp(2643) := std_logic_vector(to_signed(-25924,16));
        tmp(2644) := std_logic_vector(to_signed(-25955,16));
        tmp(2645) := std_logic_vector(to_signed(-25986,16));
        tmp(2646) := std_logic_vector(to_signed(-26016,16));
        tmp(2647) := std_logic_vector(to_signed(-26047,16));
        tmp(2648) := std_logic_vector(to_signed(-26077,16));
        tmp(2649) := std_logic_vector(to_signed(-26108,16));
        tmp(2650) := std_logic_vector(to_signed(-26138,16));
        tmp(2651) := std_logic_vector(to_signed(-26168,16));
        tmp(2652) := std_logic_vector(to_signed(-26198,16));
        tmp(2653) := std_logic_vector(to_signed(-26229,16));
        tmp(2654) := std_logic_vector(to_signed(-26259,16));
        tmp(2655) := std_logic_vector(to_signed(-26289,16));
        tmp(2656) := std_logic_vector(to_signed(-26319,16));
        tmp(2657) := std_logic_vector(to_signed(-26349,16));
        tmp(2658) := std_logic_vector(to_signed(-26378,16));
        tmp(2659) := std_logic_vector(to_signed(-26408,16));
        tmp(2660) := std_logic_vector(to_signed(-26438,16));
        tmp(2661) := std_logic_vector(to_signed(-26468,16));
        tmp(2662) := std_logic_vector(to_signed(-26497,16));
        tmp(2663) := std_logic_vector(to_signed(-26527,16));
        tmp(2664) := std_logic_vector(to_signed(-26556,16));
        tmp(2665) := std_logic_vector(to_signed(-26586,16));
        tmp(2666) := std_logic_vector(to_signed(-26615,16));
        tmp(2667) := std_logic_vector(to_signed(-26644,16));
        tmp(2668) := std_logic_vector(to_signed(-26674,16));
        tmp(2669) := std_logic_vector(to_signed(-26703,16));
        tmp(2670) := std_logic_vector(to_signed(-26732,16));
        tmp(2671) := std_logic_vector(to_signed(-26761,16));
        tmp(2672) := std_logic_vector(to_signed(-26790,16));
        tmp(2673) := std_logic_vector(to_signed(-26819,16));
        tmp(2674) := std_logic_vector(to_signed(-26848,16));
        tmp(2675) := std_logic_vector(to_signed(-26876,16));
        tmp(2676) := std_logic_vector(to_signed(-26905,16));
        tmp(2677) := std_logic_vector(to_signed(-26934,16));
        tmp(2678) := std_logic_vector(to_signed(-26962,16));
        tmp(2679) := std_logic_vector(to_signed(-26991,16));
        tmp(2680) := std_logic_vector(to_signed(-27019,16));
        tmp(2681) := std_logic_vector(to_signed(-27048,16));
        tmp(2682) := std_logic_vector(to_signed(-27076,16));
        tmp(2683) := std_logic_vector(to_signed(-27104,16));
        tmp(2684) := std_logic_vector(to_signed(-27133,16));
        tmp(2685) := std_logic_vector(to_signed(-27161,16));
        tmp(2686) := std_logic_vector(to_signed(-27189,16));
        tmp(2687) := std_logic_vector(to_signed(-27217,16));
        tmp(2688) := std_logic_vector(to_signed(-27245,16));
        tmp(2689) := std_logic_vector(to_signed(-27273,16));
        tmp(2690) := std_logic_vector(to_signed(-27300,16));
        tmp(2691) := std_logic_vector(to_signed(-27328,16));
        tmp(2692) := std_logic_vector(to_signed(-27356,16));
        tmp(2693) := std_logic_vector(to_signed(-27384,16));
        tmp(2694) := std_logic_vector(to_signed(-27411,16));
        tmp(2695) := std_logic_vector(to_signed(-27439,16));
        tmp(2696) := std_logic_vector(to_signed(-27466,16));
        tmp(2697) := std_logic_vector(to_signed(-27493,16));
        tmp(2698) := std_logic_vector(to_signed(-27521,16));
        tmp(2699) := std_logic_vector(to_signed(-27548,16));
        tmp(2700) := std_logic_vector(to_signed(-27575,16));
        tmp(2701) := std_logic_vector(to_signed(-27602,16));
        tmp(2702) := std_logic_vector(to_signed(-27629,16));
        tmp(2703) := std_logic_vector(to_signed(-27656,16));
        tmp(2704) := std_logic_vector(to_signed(-27683,16));
        tmp(2705) := std_logic_vector(to_signed(-27710,16));
        tmp(2706) := std_logic_vector(to_signed(-27737,16));
        tmp(2707) := std_logic_vector(to_signed(-27764,16));
        tmp(2708) := std_logic_vector(to_signed(-27790,16));
        tmp(2709) := std_logic_vector(to_signed(-27817,16));
        tmp(2710) := std_logic_vector(to_signed(-27843,16));
        tmp(2711) := std_logic_vector(to_signed(-27870,16));
        tmp(2712) := std_logic_vector(to_signed(-27896,16));
        tmp(2713) := std_logic_vector(to_signed(-27923,16));
        tmp(2714) := std_logic_vector(to_signed(-27949,16));
        tmp(2715) := std_logic_vector(to_signed(-27975,16));
        tmp(2716) := std_logic_vector(to_signed(-28001,16));
        tmp(2717) := std_logic_vector(to_signed(-28027,16));
        tmp(2718) := std_logic_vector(to_signed(-28053,16));
        tmp(2719) := std_logic_vector(to_signed(-28079,16));
        tmp(2720) := std_logic_vector(to_signed(-28105,16));
        tmp(2721) := std_logic_vector(to_signed(-28131,16));
        tmp(2722) := std_logic_vector(to_signed(-28157,16));
        tmp(2723) := std_logic_vector(to_signed(-28182,16));
        tmp(2724) := std_logic_vector(to_signed(-28208,16));
        tmp(2725) := std_logic_vector(to_signed(-28234,16));
        tmp(2726) := std_logic_vector(to_signed(-28259,16));
        tmp(2727) := std_logic_vector(to_signed(-28284,16));
        tmp(2728) := std_logic_vector(to_signed(-28310,16));
        tmp(2729) := std_logic_vector(to_signed(-28335,16));
        tmp(2730) := std_logic_vector(to_signed(-28360,16));
        tmp(2731) := std_logic_vector(to_signed(-28385,16));
        tmp(2732) := std_logic_vector(to_signed(-28411,16));
        tmp(2733) := std_logic_vector(to_signed(-28436,16));
        tmp(2734) := std_logic_vector(to_signed(-28460,16));
        tmp(2735) := std_logic_vector(to_signed(-28485,16));
        tmp(2736) := std_logic_vector(to_signed(-28510,16));
        tmp(2737) := std_logic_vector(to_signed(-28535,16));
        tmp(2738) := std_logic_vector(to_signed(-28560,16));
        tmp(2739) := std_logic_vector(to_signed(-28584,16));
        tmp(2740) := std_logic_vector(to_signed(-28609,16));
        tmp(2741) := std_logic_vector(to_signed(-28633,16));
        tmp(2742) := std_logic_vector(to_signed(-28658,16));
        tmp(2743) := std_logic_vector(to_signed(-28682,16));
        tmp(2744) := std_logic_vector(to_signed(-28706,16));
        tmp(2745) := std_logic_vector(to_signed(-28730,16));
        tmp(2746) := std_logic_vector(to_signed(-28755,16));
        tmp(2747) := std_logic_vector(to_signed(-28779,16));
        tmp(2748) := std_logic_vector(to_signed(-28803,16));
        tmp(2749) := std_logic_vector(to_signed(-28827,16));
        tmp(2750) := std_logic_vector(to_signed(-28850,16));
        tmp(2751) := std_logic_vector(to_signed(-28874,16));
        tmp(2752) := std_logic_vector(to_signed(-28898,16));
        tmp(2753) := std_logic_vector(to_signed(-28922,16));
        tmp(2754) := std_logic_vector(to_signed(-28945,16));
        tmp(2755) := std_logic_vector(to_signed(-28969,16));
        tmp(2756) := std_logic_vector(to_signed(-28992,16));
        tmp(2757) := std_logic_vector(to_signed(-29016,16));
        tmp(2758) := std_logic_vector(to_signed(-29039,16));
        tmp(2759) := std_logic_vector(to_signed(-29062,16));
        tmp(2760) := std_logic_vector(to_signed(-29085,16));
        tmp(2761) := std_logic_vector(to_signed(-29108,16));
        tmp(2762) := std_logic_vector(to_signed(-29131,16));
        tmp(2763) := std_logic_vector(to_signed(-29154,16));
        tmp(2764) := std_logic_vector(to_signed(-29177,16));
        tmp(2765) := std_logic_vector(to_signed(-29200,16));
        tmp(2766) := std_logic_vector(to_signed(-29223,16));
        tmp(2767) := std_logic_vector(to_signed(-29246,16));
        tmp(2768) := std_logic_vector(to_signed(-29268,16));
        tmp(2769) := std_logic_vector(to_signed(-29291,16));
        tmp(2770) := std_logic_vector(to_signed(-29313,16));
        tmp(2771) := std_logic_vector(to_signed(-29336,16));
        tmp(2772) := std_logic_vector(to_signed(-29358,16));
        tmp(2773) := std_logic_vector(to_signed(-29380,16));
        tmp(2774) := std_logic_vector(to_signed(-29403,16));
        tmp(2775) := std_logic_vector(to_signed(-29425,16));
        tmp(2776) := std_logic_vector(to_signed(-29447,16));
        tmp(2777) := std_logic_vector(to_signed(-29469,16));
        tmp(2778) := std_logic_vector(to_signed(-29491,16));
        tmp(2779) := std_logic_vector(to_signed(-29513,16));
        tmp(2780) := std_logic_vector(to_signed(-29534,16));
        tmp(2781) := std_logic_vector(to_signed(-29556,16));
        tmp(2782) := std_logic_vector(to_signed(-29578,16));
        tmp(2783) := std_logic_vector(to_signed(-29599,16));
        tmp(2784) := std_logic_vector(to_signed(-29621,16));
        tmp(2785) := std_logic_vector(to_signed(-29642,16));
        tmp(2786) := std_logic_vector(to_signed(-29664,16));
        tmp(2787) := std_logic_vector(to_signed(-29685,16));
        tmp(2788) := std_logic_vector(to_signed(-29706,16));
        tmp(2789) := std_logic_vector(to_signed(-29728,16));
        tmp(2790) := std_logic_vector(to_signed(-29749,16));
        tmp(2791) := std_logic_vector(to_signed(-29770,16));
        tmp(2792) := std_logic_vector(to_signed(-29791,16));
        tmp(2793) := std_logic_vector(to_signed(-29812,16));
        tmp(2794) := std_logic_vector(to_signed(-29832,16));
        tmp(2795) := std_logic_vector(to_signed(-29853,16));
        tmp(2796) := std_logic_vector(to_signed(-29874,16));
        tmp(2797) := std_logic_vector(to_signed(-29894,16));
        tmp(2798) := std_logic_vector(to_signed(-29915,16));
        tmp(2799) := std_logic_vector(to_signed(-29936,16));
        tmp(2800) := std_logic_vector(to_signed(-29956,16));
        tmp(2801) := std_logic_vector(to_signed(-29976,16));
        tmp(2802) := std_logic_vector(to_signed(-29997,16));
        tmp(2803) := std_logic_vector(to_signed(-30017,16));
        tmp(2804) := std_logic_vector(to_signed(-30037,16));
        tmp(2805) := std_logic_vector(to_signed(-30057,16));
        tmp(2806) := std_logic_vector(to_signed(-30077,16));
        tmp(2807) := std_logic_vector(to_signed(-30097,16));
        tmp(2808) := std_logic_vector(to_signed(-30117,16));
        tmp(2809) := std_logic_vector(to_signed(-30136,16));
        tmp(2810) := std_logic_vector(to_signed(-30156,16));
        tmp(2811) := std_logic_vector(to_signed(-30176,16));
        tmp(2812) := std_logic_vector(to_signed(-30195,16));
        tmp(2813) := std_logic_vector(to_signed(-30215,16));
        tmp(2814) := std_logic_vector(to_signed(-30234,16));
        tmp(2815) := std_logic_vector(to_signed(-30253,16));
        tmp(2816) := std_logic_vector(to_signed(-30273,16));
        tmp(2817) := std_logic_vector(to_signed(-30292,16));
        tmp(2818) := std_logic_vector(to_signed(-30311,16));
        tmp(2819) := std_logic_vector(to_signed(-30330,16));
        tmp(2820) := std_logic_vector(to_signed(-30349,16));
        tmp(2821) := std_logic_vector(to_signed(-30368,16));
        tmp(2822) := std_logic_vector(to_signed(-30387,16));
        tmp(2823) := std_logic_vector(to_signed(-30406,16));
        tmp(2824) := std_logic_vector(to_signed(-30424,16));
        tmp(2825) := std_logic_vector(to_signed(-30443,16));
        tmp(2826) := std_logic_vector(to_signed(-30462,16));
        tmp(2827) := std_logic_vector(to_signed(-30480,16));
        tmp(2828) := std_logic_vector(to_signed(-30498,16));
        tmp(2829) := std_logic_vector(to_signed(-30517,16));
        tmp(2830) := std_logic_vector(to_signed(-30535,16));
        tmp(2831) := std_logic_vector(to_signed(-30553,16));
        tmp(2832) := std_logic_vector(to_signed(-30571,16));
        tmp(2833) := std_logic_vector(to_signed(-30589,16));
        tmp(2834) := std_logic_vector(to_signed(-30607,16));
        tmp(2835) := std_logic_vector(to_signed(-30625,16));
        tmp(2836) := std_logic_vector(to_signed(-30643,16));
        tmp(2837) := std_logic_vector(to_signed(-30661,16));
        tmp(2838) := std_logic_vector(to_signed(-30679,16));
        tmp(2839) := std_logic_vector(to_signed(-30696,16));
        tmp(2840) := std_logic_vector(to_signed(-30714,16));
        tmp(2841) := std_logic_vector(to_signed(-30731,16));
        tmp(2842) := std_logic_vector(to_signed(-30749,16));
        tmp(2843) := std_logic_vector(to_signed(-30766,16));
        tmp(2844) := std_logic_vector(to_signed(-30783,16));
        tmp(2845) := std_logic_vector(to_signed(-30800,16));
        tmp(2846) := std_logic_vector(to_signed(-30818,16));
        tmp(2847) := std_logic_vector(to_signed(-30835,16));
        tmp(2848) := std_logic_vector(to_signed(-30852,16));
        tmp(2849) := std_logic_vector(to_signed(-30868,16));
        tmp(2850) := std_logic_vector(to_signed(-30885,16));
        tmp(2851) := std_logic_vector(to_signed(-30902,16));
        tmp(2852) := std_logic_vector(to_signed(-30919,16));
        tmp(2853) := std_logic_vector(to_signed(-30935,16));
        tmp(2854) := std_logic_vector(to_signed(-30952,16));
        tmp(2855) := std_logic_vector(to_signed(-30968,16));
        tmp(2856) := std_logic_vector(to_signed(-30985,16));
        tmp(2857) := std_logic_vector(to_signed(-31001,16));
        tmp(2858) := std_logic_vector(to_signed(-31017,16));
        tmp(2859) := std_logic_vector(to_signed(-31033,16));
        tmp(2860) := std_logic_vector(to_signed(-31050,16));
        tmp(2861) := std_logic_vector(to_signed(-31066,16));
        tmp(2862) := std_logic_vector(to_signed(-31082,16));
        tmp(2863) := std_logic_vector(to_signed(-31097,16));
        tmp(2864) := std_logic_vector(to_signed(-31113,16));
        tmp(2865) := std_logic_vector(to_signed(-31129,16));
        tmp(2866) := std_logic_vector(to_signed(-31145,16));
        tmp(2867) := std_logic_vector(to_signed(-31160,16));
        tmp(2868) := std_logic_vector(to_signed(-31176,16));
        tmp(2869) := std_logic_vector(to_signed(-31191,16));
        tmp(2870) := std_logic_vector(to_signed(-31206,16));
        tmp(2871) := std_logic_vector(to_signed(-31222,16));
        tmp(2872) := std_logic_vector(to_signed(-31237,16));
        tmp(2873) := std_logic_vector(to_signed(-31252,16));
        tmp(2874) := std_logic_vector(to_signed(-31267,16));
        tmp(2875) := std_logic_vector(to_signed(-31282,16));
        tmp(2876) := std_logic_vector(to_signed(-31297,16));
        tmp(2877) := std_logic_vector(to_signed(-31312,16));
        tmp(2878) := std_logic_vector(to_signed(-31327,16));
        tmp(2879) := std_logic_vector(to_signed(-31341,16));
        tmp(2880) := std_logic_vector(to_signed(-31356,16));
        tmp(2881) := std_logic_vector(to_signed(-31371,16));
        tmp(2882) := std_logic_vector(to_signed(-31385,16));
        tmp(2883) := std_logic_vector(to_signed(-31400,16));
        tmp(2884) := std_logic_vector(to_signed(-31414,16));
        tmp(2885) := std_logic_vector(to_signed(-31428,16));
        tmp(2886) := std_logic_vector(to_signed(-31442,16));
        tmp(2887) := std_logic_vector(to_signed(-31456,16));
        tmp(2888) := std_logic_vector(to_signed(-31470,16));
        tmp(2889) := std_logic_vector(to_signed(-31484,16));
        tmp(2890) := std_logic_vector(to_signed(-31498,16));
        tmp(2891) := std_logic_vector(to_signed(-31512,16));
        tmp(2892) := std_logic_vector(to_signed(-31526,16));
        tmp(2893) := std_logic_vector(to_signed(-31539,16));
        tmp(2894) := std_logic_vector(to_signed(-31553,16));
        tmp(2895) := std_logic_vector(to_signed(-31567,16));
        tmp(2896) := std_logic_vector(to_signed(-31580,16));
        tmp(2897) := std_logic_vector(to_signed(-31593,16));
        tmp(2898) := std_logic_vector(to_signed(-31607,16));
        tmp(2899) := std_logic_vector(to_signed(-31620,16));
        tmp(2900) := std_logic_vector(to_signed(-31633,16));
        tmp(2901) := std_logic_vector(to_signed(-31646,16));
        tmp(2902) := std_logic_vector(to_signed(-31659,16));
        tmp(2903) := std_logic_vector(to_signed(-31672,16));
        tmp(2904) := std_logic_vector(to_signed(-31685,16));
        tmp(2905) := std_logic_vector(to_signed(-31698,16));
        tmp(2906) := std_logic_vector(to_signed(-31710,16));
        tmp(2907) := std_logic_vector(to_signed(-31723,16));
        tmp(2908) := std_logic_vector(to_signed(-31736,16));
        tmp(2909) := std_logic_vector(to_signed(-31748,16));
        tmp(2910) := std_logic_vector(to_signed(-31760,16));
        tmp(2911) := std_logic_vector(to_signed(-31773,16));
        tmp(2912) := std_logic_vector(to_signed(-31785,16));
        tmp(2913) := std_logic_vector(to_signed(-31797,16));
        tmp(2914) := std_logic_vector(to_signed(-31809,16));
        tmp(2915) := std_logic_vector(to_signed(-31821,16));
        tmp(2916) := std_logic_vector(to_signed(-31833,16));
        tmp(2917) := std_logic_vector(to_signed(-31845,16));
        tmp(2918) := std_logic_vector(to_signed(-31857,16));
        tmp(2919) := std_logic_vector(to_signed(-31869,16));
        tmp(2920) := std_logic_vector(to_signed(-31880,16));
        tmp(2921) := std_logic_vector(to_signed(-31892,16));
        tmp(2922) := std_logic_vector(to_signed(-31903,16));
        tmp(2923) := std_logic_vector(to_signed(-31915,16));
        tmp(2924) := std_logic_vector(to_signed(-31926,16));
        tmp(2925) := std_logic_vector(to_signed(-31937,16));
        tmp(2926) := std_logic_vector(to_signed(-31949,16));
        tmp(2927) := std_logic_vector(to_signed(-31960,16));
        tmp(2928) := std_logic_vector(to_signed(-31971,16));
        tmp(2929) := std_logic_vector(to_signed(-31982,16));
        tmp(2930) := std_logic_vector(to_signed(-31993,16));
        tmp(2931) := std_logic_vector(to_signed(-32004,16));
        tmp(2932) := std_logic_vector(to_signed(-32014,16));
        tmp(2933) := std_logic_vector(to_signed(-32025,16));
        tmp(2934) := std_logic_vector(to_signed(-32036,16));
        tmp(2935) := std_logic_vector(to_signed(-32046,16));
        tmp(2936) := std_logic_vector(to_signed(-32057,16));
        tmp(2937) := std_logic_vector(to_signed(-32067,16));
        tmp(2938) := std_logic_vector(to_signed(-32077,16));
        tmp(2939) := std_logic_vector(to_signed(-32087,16));
        tmp(2940) := std_logic_vector(to_signed(-32098,16));
        tmp(2941) := std_logic_vector(to_signed(-32108,16));
        tmp(2942) := std_logic_vector(to_signed(-32118,16));
        tmp(2943) := std_logic_vector(to_signed(-32128,16));
        tmp(2944) := std_logic_vector(to_signed(-32137,16));
        tmp(2945) := std_logic_vector(to_signed(-32147,16));
        tmp(2946) := std_logic_vector(to_signed(-32157,16));
        tmp(2947) := std_logic_vector(to_signed(-32166,16));
        tmp(2948) := std_logic_vector(to_signed(-32176,16));
        tmp(2949) := std_logic_vector(to_signed(-32185,16));
        tmp(2950) := std_logic_vector(to_signed(-32195,16));
        tmp(2951) := std_logic_vector(to_signed(-32204,16));
        tmp(2952) := std_logic_vector(to_signed(-32213,16));
        tmp(2953) := std_logic_vector(to_signed(-32223,16));
        tmp(2954) := std_logic_vector(to_signed(-32232,16));
        tmp(2955) := std_logic_vector(to_signed(-32241,16));
        tmp(2956) := std_logic_vector(to_signed(-32250,16));
        tmp(2957) := std_logic_vector(to_signed(-32258,16));
        tmp(2958) := std_logic_vector(to_signed(-32267,16));
        tmp(2959) := std_logic_vector(to_signed(-32276,16));
        tmp(2960) := std_logic_vector(to_signed(-32285,16));
        tmp(2961) := std_logic_vector(to_signed(-32293,16));
        tmp(2962) := std_logic_vector(to_signed(-32302,16));
        tmp(2963) := std_logic_vector(to_signed(-32310,16));
        tmp(2964) := std_logic_vector(to_signed(-32318,16));
        tmp(2965) := std_logic_vector(to_signed(-32327,16));
        tmp(2966) := std_logic_vector(to_signed(-32335,16));
        tmp(2967) := std_logic_vector(to_signed(-32343,16));
        tmp(2968) := std_logic_vector(to_signed(-32351,16));
        tmp(2969) := std_logic_vector(to_signed(-32359,16));
        tmp(2970) := std_logic_vector(to_signed(-32367,16));
        tmp(2971) := std_logic_vector(to_signed(-32375,16));
        tmp(2972) := std_logic_vector(to_signed(-32382,16));
        tmp(2973) := std_logic_vector(to_signed(-32390,16));
        tmp(2974) := std_logic_vector(to_signed(-32397,16));
        tmp(2975) := std_logic_vector(to_signed(-32405,16));
        tmp(2976) := std_logic_vector(to_signed(-32412,16));
        tmp(2977) := std_logic_vector(to_signed(-32420,16));
        tmp(2978) := std_logic_vector(to_signed(-32427,16));
        tmp(2979) := std_logic_vector(to_signed(-32434,16));
        tmp(2980) := std_logic_vector(to_signed(-32441,16));
        tmp(2981) := std_logic_vector(to_signed(-32448,16));
        tmp(2982) := std_logic_vector(to_signed(-32455,16));
        tmp(2983) := std_logic_vector(to_signed(-32462,16));
        tmp(2984) := std_logic_vector(to_signed(-32469,16));
        tmp(2985) := std_logic_vector(to_signed(-32476,16));
        tmp(2986) := std_logic_vector(to_signed(-32482,16));
        tmp(2987) := std_logic_vector(to_signed(-32489,16));
        tmp(2988) := std_logic_vector(to_signed(-32495,16));
        tmp(2989) := std_logic_vector(to_signed(-32502,16));
        tmp(2990) := std_logic_vector(to_signed(-32508,16));
        tmp(2991) := std_logic_vector(to_signed(-32514,16));
        tmp(2992) := std_logic_vector(to_signed(-32521,16));
        tmp(2993) := std_logic_vector(to_signed(-32527,16));
        tmp(2994) := std_logic_vector(to_signed(-32533,16));
        tmp(2995) := std_logic_vector(to_signed(-32539,16));
        tmp(2996) := std_logic_vector(to_signed(-32545,16));
        tmp(2997) := std_logic_vector(to_signed(-32550,16));
        tmp(2998) := std_logic_vector(to_signed(-32556,16));
        tmp(2999) := std_logic_vector(to_signed(-32562,16));
        tmp(3000) := std_logic_vector(to_signed(-32567,16));
        tmp(3001) := std_logic_vector(to_signed(-32573,16));
        tmp(3002) := std_logic_vector(to_signed(-32578,16));
        tmp(3003) := std_logic_vector(to_signed(-32584,16));
        tmp(3004) := std_logic_vector(to_signed(-32589,16));
        tmp(3005) := std_logic_vector(to_signed(-32594,16));
        tmp(3006) := std_logic_vector(to_signed(-32599,16));
        tmp(3007) := std_logic_vector(to_signed(-32604,16));
        tmp(3008) := std_logic_vector(to_signed(-32609,16));
        tmp(3009) := std_logic_vector(to_signed(-32614,16));
        tmp(3010) := std_logic_vector(to_signed(-32619,16));
        tmp(3011) := std_logic_vector(to_signed(-32624,16));
        tmp(3012) := std_logic_vector(to_signed(-32628,16));
        tmp(3013) := std_logic_vector(to_signed(-32633,16));
        tmp(3014) := std_logic_vector(to_signed(-32637,16));
        tmp(3015) := std_logic_vector(to_signed(-32642,16));
        tmp(3016) := std_logic_vector(to_signed(-32646,16));
        tmp(3017) := std_logic_vector(to_signed(-32650,16));
        tmp(3018) := std_logic_vector(to_signed(-32655,16));
        tmp(3019) := std_logic_vector(to_signed(-32659,16));
        tmp(3020) := std_logic_vector(to_signed(-32663,16));
        tmp(3021) := std_logic_vector(to_signed(-32667,16));
        tmp(3022) := std_logic_vector(to_signed(-32671,16));
        tmp(3023) := std_logic_vector(to_signed(-32674,16));
        tmp(3024) := std_logic_vector(to_signed(-32678,16));
        tmp(3025) := std_logic_vector(to_signed(-32682,16));
        tmp(3026) := std_logic_vector(to_signed(-32685,16));
        tmp(3027) := std_logic_vector(to_signed(-32689,16));
        tmp(3028) := std_logic_vector(to_signed(-32692,16));
        tmp(3029) := std_logic_vector(to_signed(-32696,16));
        tmp(3030) := std_logic_vector(to_signed(-32699,16));
        tmp(3031) := std_logic_vector(to_signed(-32702,16));
        tmp(3032) := std_logic_vector(to_signed(-32705,16));
        tmp(3033) := std_logic_vector(to_signed(-32708,16));
        tmp(3034) := std_logic_vector(to_signed(-32711,16));
        tmp(3035) := std_logic_vector(to_signed(-32714,16));
        tmp(3036) := std_logic_vector(to_signed(-32717,16));
        tmp(3037) := std_logic_vector(to_signed(-32720,16));
        tmp(3038) := std_logic_vector(to_signed(-32722,16));
        tmp(3039) := std_logic_vector(to_signed(-32725,16));
        tmp(3040) := std_logic_vector(to_signed(-32728,16));
        tmp(3041) := std_logic_vector(to_signed(-32730,16));
        tmp(3042) := std_logic_vector(to_signed(-32732,16));
        tmp(3043) := std_logic_vector(to_signed(-32735,16));
        tmp(3044) := std_logic_vector(to_signed(-32737,16));
        tmp(3045) := std_logic_vector(to_signed(-32739,16));
        tmp(3046) := std_logic_vector(to_signed(-32741,16));
        tmp(3047) := std_logic_vector(to_signed(-32743,16));
        tmp(3048) := std_logic_vector(to_signed(-32745,16));
        tmp(3049) := std_logic_vector(to_signed(-32747,16));
        tmp(3050) := std_logic_vector(to_signed(-32748,16));
        tmp(3051) := std_logic_vector(to_signed(-32750,16));
        tmp(3052) := std_logic_vector(to_signed(-32752,16));
        tmp(3053) := std_logic_vector(to_signed(-32753,16));
        tmp(3054) := std_logic_vector(to_signed(-32755,16));
        tmp(3055) := std_logic_vector(to_signed(-32756,16));
        tmp(3056) := std_logic_vector(to_signed(-32757,16));
        tmp(3057) := std_logic_vector(to_signed(-32758,16));
        tmp(3058) := std_logic_vector(to_signed(-32759,16));
        tmp(3059) := std_logic_vector(to_signed(-32760,16));
        tmp(3060) := std_logic_vector(to_signed(-32761,16));
        tmp(3061) := std_logic_vector(to_signed(-32762,16));
        tmp(3062) := std_logic_vector(to_signed(-32763,16));
        tmp(3063) := std_logic_vector(to_signed(-32764,16));
        tmp(3064) := std_logic_vector(to_signed(-32765,16));
        tmp(3065) := std_logic_vector(to_signed(-32765,16));
        tmp(3066) := std_logic_vector(to_signed(-32766,16));
        tmp(3067) := std_logic_vector(to_signed(-32766,16));
        tmp(3068) := std_logic_vector(to_signed(-32766,16));
        tmp(3069) := std_logic_vector(to_signed(-32767,16));
        tmp(3070) := std_logic_vector(to_signed(-32767,16));
        tmp(3071) := std_logic_vector(to_signed(-32767,16));
        tmp(3072) := std_logic_vector(to_signed(-32767,16));
        tmp(3073) := std_logic_vector(to_signed(-32767,16));
        tmp(3074) := std_logic_vector(to_signed(-32767,16));
        tmp(3075) := std_logic_vector(to_signed(-32767,16));
        tmp(3076) := std_logic_vector(to_signed(-32766,16));
        tmp(3077) := std_logic_vector(to_signed(-32766,16));
        tmp(3078) := std_logic_vector(to_signed(-32766,16));
        tmp(3079) := std_logic_vector(to_signed(-32765,16));
        tmp(3080) := std_logic_vector(to_signed(-32765,16));
        tmp(3081) := std_logic_vector(to_signed(-32764,16));
        tmp(3082) := std_logic_vector(to_signed(-32763,16));
        tmp(3083) := std_logic_vector(to_signed(-32762,16));
        tmp(3084) := std_logic_vector(to_signed(-32761,16));
        tmp(3085) := std_logic_vector(to_signed(-32760,16));
        tmp(3086) := std_logic_vector(to_signed(-32759,16));
        tmp(3087) := std_logic_vector(to_signed(-32758,16));
        tmp(3088) := std_logic_vector(to_signed(-32757,16));
        tmp(3089) := std_logic_vector(to_signed(-32756,16));
        tmp(3090) := std_logic_vector(to_signed(-32755,16));
        tmp(3091) := std_logic_vector(to_signed(-32753,16));
        tmp(3092) := std_logic_vector(to_signed(-32752,16));
        tmp(3093) := std_logic_vector(to_signed(-32750,16));
        tmp(3094) := std_logic_vector(to_signed(-32748,16));
        tmp(3095) := std_logic_vector(to_signed(-32747,16));
        tmp(3096) := std_logic_vector(to_signed(-32745,16));
        tmp(3097) := std_logic_vector(to_signed(-32743,16));
        tmp(3098) := std_logic_vector(to_signed(-32741,16));
        tmp(3099) := std_logic_vector(to_signed(-32739,16));
        tmp(3100) := std_logic_vector(to_signed(-32737,16));
        tmp(3101) := std_logic_vector(to_signed(-32735,16));
        tmp(3102) := std_logic_vector(to_signed(-32732,16));
        tmp(3103) := std_logic_vector(to_signed(-32730,16));
        tmp(3104) := std_logic_vector(to_signed(-32728,16));
        tmp(3105) := std_logic_vector(to_signed(-32725,16));
        tmp(3106) := std_logic_vector(to_signed(-32722,16));
        tmp(3107) := std_logic_vector(to_signed(-32720,16));
        tmp(3108) := std_logic_vector(to_signed(-32717,16));
        tmp(3109) := std_logic_vector(to_signed(-32714,16));
        tmp(3110) := std_logic_vector(to_signed(-32711,16));
        tmp(3111) := std_logic_vector(to_signed(-32708,16));
        tmp(3112) := std_logic_vector(to_signed(-32705,16));
        tmp(3113) := std_logic_vector(to_signed(-32702,16));
        tmp(3114) := std_logic_vector(to_signed(-32699,16));
        tmp(3115) := std_logic_vector(to_signed(-32696,16));
        tmp(3116) := std_logic_vector(to_signed(-32692,16));
        tmp(3117) := std_logic_vector(to_signed(-32689,16));
        tmp(3118) := std_logic_vector(to_signed(-32685,16));
        tmp(3119) := std_logic_vector(to_signed(-32682,16));
        tmp(3120) := std_logic_vector(to_signed(-32678,16));
        tmp(3121) := std_logic_vector(to_signed(-32674,16));
        tmp(3122) := std_logic_vector(to_signed(-32671,16));
        tmp(3123) := std_logic_vector(to_signed(-32667,16));
        tmp(3124) := std_logic_vector(to_signed(-32663,16));
        tmp(3125) := std_logic_vector(to_signed(-32659,16));
        tmp(3126) := std_logic_vector(to_signed(-32655,16));
        tmp(3127) := std_logic_vector(to_signed(-32650,16));
        tmp(3128) := std_logic_vector(to_signed(-32646,16));
        tmp(3129) := std_logic_vector(to_signed(-32642,16));
        tmp(3130) := std_logic_vector(to_signed(-32637,16));
        tmp(3131) := std_logic_vector(to_signed(-32633,16));
        tmp(3132) := std_logic_vector(to_signed(-32628,16));
        tmp(3133) := std_logic_vector(to_signed(-32624,16));
        tmp(3134) := std_logic_vector(to_signed(-32619,16));
        tmp(3135) := std_logic_vector(to_signed(-32614,16));
        tmp(3136) := std_logic_vector(to_signed(-32609,16));
        tmp(3137) := std_logic_vector(to_signed(-32604,16));
        tmp(3138) := std_logic_vector(to_signed(-32599,16));
        tmp(3139) := std_logic_vector(to_signed(-32594,16));
        tmp(3140) := std_logic_vector(to_signed(-32589,16));
        tmp(3141) := std_logic_vector(to_signed(-32584,16));
        tmp(3142) := std_logic_vector(to_signed(-32578,16));
        tmp(3143) := std_logic_vector(to_signed(-32573,16));
        tmp(3144) := std_logic_vector(to_signed(-32567,16));
        tmp(3145) := std_logic_vector(to_signed(-32562,16));
        tmp(3146) := std_logic_vector(to_signed(-32556,16));
        tmp(3147) := std_logic_vector(to_signed(-32550,16));
        tmp(3148) := std_logic_vector(to_signed(-32545,16));
        tmp(3149) := std_logic_vector(to_signed(-32539,16));
        tmp(3150) := std_logic_vector(to_signed(-32533,16));
        tmp(3151) := std_logic_vector(to_signed(-32527,16));
        tmp(3152) := std_logic_vector(to_signed(-32521,16));
        tmp(3153) := std_logic_vector(to_signed(-32514,16));
        tmp(3154) := std_logic_vector(to_signed(-32508,16));
        tmp(3155) := std_logic_vector(to_signed(-32502,16));
        tmp(3156) := std_logic_vector(to_signed(-32495,16));
        tmp(3157) := std_logic_vector(to_signed(-32489,16));
        tmp(3158) := std_logic_vector(to_signed(-32482,16));
        tmp(3159) := std_logic_vector(to_signed(-32476,16));
        tmp(3160) := std_logic_vector(to_signed(-32469,16));
        tmp(3161) := std_logic_vector(to_signed(-32462,16));
        tmp(3162) := std_logic_vector(to_signed(-32455,16));
        tmp(3163) := std_logic_vector(to_signed(-32448,16));
        tmp(3164) := std_logic_vector(to_signed(-32441,16));
        tmp(3165) := std_logic_vector(to_signed(-32434,16));
        tmp(3166) := std_logic_vector(to_signed(-32427,16));
        tmp(3167) := std_logic_vector(to_signed(-32420,16));
        tmp(3168) := std_logic_vector(to_signed(-32412,16));
        tmp(3169) := std_logic_vector(to_signed(-32405,16));
        tmp(3170) := std_logic_vector(to_signed(-32397,16));
        tmp(3171) := std_logic_vector(to_signed(-32390,16));
        tmp(3172) := std_logic_vector(to_signed(-32382,16));
        tmp(3173) := std_logic_vector(to_signed(-32375,16));
        tmp(3174) := std_logic_vector(to_signed(-32367,16));
        tmp(3175) := std_logic_vector(to_signed(-32359,16));
        tmp(3176) := std_logic_vector(to_signed(-32351,16));
        tmp(3177) := std_logic_vector(to_signed(-32343,16));
        tmp(3178) := std_logic_vector(to_signed(-32335,16));
        tmp(3179) := std_logic_vector(to_signed(-32327,16));
        tmp(3180) := std_logic_vector(to_signed(-32318,16));
        tmp(3181) := std_logic_vector(to_signed(-32310,16));
        tmp(3182) := std_logic_vector(to_signed(-32302,16));
        tmp(3183) := std_logic_vector(to_signed(-32293,16));
        tmp(3184) := std_logic_vector(to_signed(-32285,16));
        tmp(3185) := std_logic_vector(to_signed(-32276,16));
        tmp(3186) := std_logic_vector(to_signed(-32267,16));
        tmp(3187) := std_logic_vector(to_signed(-32258,16));
        tmp(3188) := std_logic_vector(to_signed(-32250,16));
        tmp(3189) := std_logic_vector(to_signed(-32241,16));
        tmp(3190) := std_logic_vector(to_signed(-32232,16));
        tmp(3191) := std_logic_vector(to_signed(-32223,16));
        tmp(3192) := std_logic_vector(to_signed(-32213,16));
        tmp(3193) := std_logic_vector(to_signed(-32204,16));
        tmp(3194) := std_logic_vector(to_signed(-32195,16));
        tmp(3195) := std_logic_vector(to_signed(-32185,16));
        tmp(3196) := std_logic_vector(to_signed(-32176,16));
        tmp(3197) := std_logic_vector(to_signed(-32166,16));
        tmp(3198) := std_logic_vector(to_signed(-32157,16));
        tmp(3199) := std_logic_vector(to_signed(-32147,16));
        tmp(3200) := std_logic_vector(to_signed(-32137,16));
        tmp(3201) := std_logic_vector(to_signed(-32128,16));
        tmp(3202) := std_logic_vector(to_signed(-32118,16));
        tmp(3203) := std_logic_vector(to_signed(-32108,16));
        tmp(3204) := std_logic_vector(to_signed(-32098,16));
        tmp(3205) := std_logic_vector(to_signed(-32087,16));
        tmp(3206) := std_logic_vector(to_signed(-32077,16));
        tmp(3207) := std_logic_vector(to_signed(-32067,16));
        tmp(3208) := std_logic_vector(to_signed(-32057,16));
        tmp(3209) := std_logic_vector(to_signed(-32046,16));
        tmp(3210) := std_logic_vector(to_signed(-32036,16));
        tmp(3211) := std_logic_vector(to_signed(-32025,16));
        tmp(3212) := std_logic_vector(to_signed(-32014,16));
        tmp(3213) := std_logic_vector(to_signed(-32004,16));
        tmp(3214) := std_logic_vector(to_signed(-31993,16));
        tmp(3215) := std_logic_vector(to_signed(-31982,16));
        tmp(3216) := std_logic_vector(to_signed(-31971,16));
        tmp(3217) := std_logic_vector(to_signed(-31960,16));
        tmp(3218) := std_logic_vector(to_signed(-31949,16));
        tmp(3219) := std_logic_vector(to_signed(-31937,16));
        tmp(3220) := std_logic_vector(to_signed(-31926,16));
        tmp(3221) := std_logic_vector(to_signed(-31915,16));
        tmp(3222) := std_logic_vector(to_signed(-31903,16));
        tmp(3223) := std_logic_vector(to_signed(-31892,16));
        tmp(3224) := std_logic_vector(to_signed(-31880,16));
        tmp(3225) := std_logic_vector(to_signed(-31869,16));
        tmp(3226) := std_logic_vector(to_signed(-31857,16));
        tmp(3227) := std_logic_vector(to_signed(-31845,16));
        tmp(3228) := std_logic_vector(to_signed(-31833,16));
        tmp(3229) := std_logic_vector(to_signed(-31821,16));
        tmp(3230) := std_logic_vector(to_signed(-31809,16));
        tmp(3231) := std_logic_vector(to_signed(-31797,16));
        tmp(3232) := std_logic_vector(to_signed(-31785,16));
        tmp(3233) := std_logic_vector(to_signed(-31773,16));
        tmp(3234) := std_logic_vector(to_signed(-31760,16));
        tmp(3235) := std_logic_vector(to_signed(-31748,16));
        tmp(3236) := std_logic_vector(to_signed(-31736,16));
        tmp(3237) := std_logic_vector(to_signed(-31723,16));
        tmp(3238) := std_logic_vector(to_signed(-31710,16));
        tmp(3239) := std_logic_vector(to_signed(-31698,16));
        tmp(3240) := std_logic_vector(to_signed(-31685,16));
        tmp(3241) := std_logic_vector(to_signed(-31672,16));
        tmp(3242) := std_logic_vector(to_signed(-31659,16));
        tmp(3243) := std_logic_vector(to_signed(-31646,16));
        tmp(3244) := std_logic_vector(to_signed(-31633,16));
        tmp(3245) := std_logic_vector(to_signed(-31620,16));
        tmp(3246) := std_logic_vector(to_signed(-31607,16));
        tmp(3247) := std_logic_vector(to_signed(-31593,16));
        tmp(3248) := std_logic_vector(to_signed(-31580,16));
        tmp(3249) := std_logic_vector(to_signed(-31567,16));
        tmp(3250) := std_logic_vector(to_signed(-31553,16));
        tmp(3251) := std_logic_vector(to_signed(-31539,16));
        tmp(3252) := std_logic_vector(to_signed(-31526,16));
        tmp(3253) := std_logic_vector(to_signed(-31512,16));
        tmp(3254) := std_logic_vector(to_signed(-31498,16));
        tmp(3255) := std_logic_vector(to_signed(-31484,16));
        tmp(3256) := std_logic_vector(to_signed(-31470,16));
        tmp(3257) := std_logic_vector(to_signed(-31456,16));
        tmp(3258) := std_logic_vector(to_signed(-31442,16));
        tmp(3259) := std_logic_vector(to_signed(-31428,16));
        tmp(3260) := std_logic_vector(to_signed(-31414,16));
        tmp(3261) := std_logic_vector(to_signed(-31400,16));
        tmp(3262) := std_logic_vector(to_signed(-31385,16));
        tmp(3263) := std_logic_vector(to_signed(-31371,16));
        tmp(3264) := std_logic_vector(to_signed(-31356,16));
        tmp(3265) := std_logic_vector(to_signed(-31341,16));
        tmp(3266) := std_logic_vector(to_signed(-31327,16));
        tmp(3267) := std_logic_vector(to_signed(-31312,16));
        tmp(3268) := std_logic_vector(to_signed(-31297,16));
        tmp(3269) := std_logic_vector(to_signed(-31282,16));
        tmp(3270) := std_logic_vector(to_signed(-31267,16));
        tmp(3271) := std_logic_vector(to_signed(-31252,16));
        tmp(3272) := std_logic_vector(to_signed(-31237,16));
        tmp(3273) := std_logic_vector(to_signed(-31222,16));
        tmp(3274) := std_logic_vector(to_signed(-31206,16));
        tmp(3275) := std_logic_vector(to_signed(-31191,16));
        tmp(3276) := std_logic_vector(to_signed(-31176,16));
        tmp(3277) := std_logic_vector(to_signed(-31160,16));
        tmp(3278) := std_logic_vector(to_signed(-31145,16));
        tmp(3279) := std_logic_vector(to_signed(-31129,16));
        tmp(3280) := std_logic_vector(to_signed(-31113,16));
        tmp(3281) := std_logic_vector(to_signed(-31097,16));
        tmp(3282) := std_logic_vector(to_signed(-31082,16));
        tmp(3283) := std_logic_vector(to_signed(-31066,16));
        tmp(3284) := std_logic_vector(to_signed(-31050,16));
        tmp(3285) := std_logic_vector(to_signed(-31033,16));
        tmp(3286) := std_logic_vector(to_signed(-31017,16));
        tmp(3287) := std_logic_vector(to_signed(-31001,16));
        tmp(3288) := std_logic_vector(to_signed(-30985,16));
        tmp(3289) := std_logic_vector(to_signed(-30968,16));
        tmp(3290) := std_logic_vector(to_signed(-30952,16));
        tmp(3291) := std_logic_vector(to_signed(-30935,16));
        tmp(3292) := std_logic_vector(to_signed(-30919,16));
        tmp(3293) := std_logic_vector(to_signed(-30902,16));
        tmp(3294) := std_logic_vector(to_signed(-30885,16));
        tmp(3295) := std_logic_vector(to_signed(-30868,16));
        tmp(3296) := std_logic_vector(to_signed(-30852,16));
        tmp(3297) := std_logic_vector(to_signed(-30835,16));
        tmp(3298) := std_logic_vector(to_signed(-30818,16));
        tmp(3299) := std_logic_vector(to_signed(-30800,16));
        tmp(3300) := std_logic_vector(to_signed(-30783,16));
        tmp(3301) := std_logic_vector(to_signed(-30766,16));
        tmp(3302) := std_logic_vector(to_signed(-30749,16));
        tmp(3303) := std_logic_vector(to_signed(-30731,16));
        tmp(3304) := std_logic_vector(to_signed(-30714,16));
        tmp(3305) := std_logic_vector(to_signed(-30696,16));
        tmp(3306) := std_logic_vector(to_signed(-30679,16));
        tmp(3307) := std_logic_vector(to_signed(-30661,16));
        tmp(3308) := std_logic_vector(to_signed(-30643,16));
        tmp(3309) := std_logic_vector(to_signed(-30625,16));
        tmp(3310) := std_logic_vector(to_signed(-30607,16));
        tmp(3311) := std_logic_vector(to_signed(-30589,16));
        tmp(3312) := std_logic_vector(to_signed(-30571,16));
        tmp(3313) := std_logic_vector(to_signed(-30553,16));
        tmp(3314) := std_logic_vector(to_signed(-30535,16));
        tmp(3315) := std_logic_vector(to_signed(-30517,16));
        tmp(3316) := std_logic_vector(to_signed(-30498,16));
        tmp(3317) := std_logic_vector(to_signed(-30480,16));
        tmp(3318) := std_logic_vector(to_signed(-30462,16));
        tmp(3319) := std_logic_vector(to_signed(-30443,16));
        tmp(3320) := std_logic_vector(to_signed(-30424,16));
        tmp(3321) := std_logic_vector(to_signed(-30406,16));
        tmp(3322) := std_logic_vector(to_signed(-30387,16));
        tmp(3323) := std_logic_vector(to_signed(-30368,16));
        tmp(3324) := std_logic_vector(to_signed(-30349,16));
        tmp(3325) := std_logic_vector(to_signed(-30330,16));
        tmp(3326) := std_logic_vector(to_signed(-30311,16));
        tmp(3327) := std_logic_vector(to_signed(-30292,16));
        tmp(3328) := std_logic_vector(to_signed(-30273,16));
        tmp(3329) := std_logic_vector(to_signed(-30253,16));
        tmp(3330) := std_logic_vector(to_signed(-30234,16));
        tmp(3331) := std_logic_vector(to_signed(-30215,16));
        tmp(3332) := std_logic_vector(to_signed(-30195,16));
        tmp(3333) := std_logic_vector(to_signed(-30176,16));
        tmp(3334) := std_logic_vector(to_signed(-30156,16));
        tmp(3335) := std_logic_vector(to_signed(-30136,16));
        tmp(3336) := std_logic_vector(to_signed(-30117,16));
        tmp(3337) := std_logic_vector(to_signed(-30097,16));
        tmp(3338) := std_logic_vector(to_signed(-30077,16));
        tmp(3339) := std_logic_vector(to_signed(-30057,16));
        tmp(3340) := std_logic_vector(to_signed(-30037,16));
        tmp(3341) := std_logic_vector(to_signed(-30017,16));
        tmp(3342) := std_logic_vector(to_signed(-29997,16));
        tmp(3343) := std_logic_vector(to_signed(-29976,16));
        tmp(3344) := std_logic_vector(to_signed(-29956,16));
        tmp(3345) := std_logic_vector(to_signed(-29936,16));
        tmp(3346) := std_logic_vector(to_signed(-29915,16));
        tmp(3347) := std_logic_vector(to_signed(-29894,16));
        tmp(3348) := std_logic_vector(to_signed(-29874,16));
        tmp(3349) := std_logic_vector(to_signed(-29853,16));
        tmp(3350) := std_logic_vector(to_signed(-29832,16));
        tmp(3351) := std_logic_vector(to_signed(-29812,16));
        tmp(3352) := std_logic_vector(to_signed(-29791,16));
        tmp(3353) := std_logic_vector(to_signed(-29770,16));
        tmp(3354) := std_logic_vector(to_signed(-29749,16));
        tmp(3355) := std_logic_vector(to_signed(-29728,16));
        tmp(3356) := std_logic_vector(to_signed(-29706,16));
        tmp(3357) := std_logic_vector(to_signed(-29685,16));
        tmp(3358) := std_logic_vector(to_signed(-29664,16));
        tmp(3359) := std_logic_vector(to_signed(-29642,16));
        tmp(3360) := std_logic_vector(to_signed(-29621,16));
        tmp(3361) := std_logic_vector(to_signed(-29599,16));
        tmp(3362) := std_logic_vector(to_signed(-29578,16));
        tmp(3363) := std_logic_vector(to_signed(-29556,16));
        tmp(3364) := std_logic_vector(to_signed(-29534,16));
        tmp(3365) := std_logic_vector(to_signed(-29513,16));
        tmp(3366) := std_logic_vector(to_signed(-29491,16));
        tmp(3367) := std_logic_vector(to_signed(-29469,16));
        tmp(3368) := std_logic_vector(to_signed(-29447,16));
        tmp(3369) := std_logic_vector(to_signed(-29425,16));
        tmp(3370) := std_logic_vector(to_signed(-29403,16));
        tmp(3371) := std_logic_vector(to_signed(-29380,16));
        tmp(3372) := std_logic_vector(to_signed(-29358,16));
        tmp(3373) := std_logic_vector(to_signed(-29336,16));
        tmp(3374) := std_logic_vector(to_signed(-29313,16));
        tmp(3375) := std_logic_vector(to_signed(-29291,16));
        tmp(3376) := std_logic_vector(to_signed(-29268,16));
        tmp(3377) := std_logic_vector(to_signed(-29246,16));
        tmp(3378) := std_logic_vector(to_signed(-29223,16));
        tmp(3379) := std_logic_vector(to_signed(-29200,16));
        tmp(3380) := std_logic_vector(to_signed(-29177,16));
        tmp(3381) := std_logic_vector(to_signed(-29154,16));
        tmp(3382) := std_logic_vector(to_signed(-29131,16));
        tmp(3383) := std_logic_vector(to_signed(-29108,16));
        tmp(3384) := std_logic_vector(to_signed(-29085,16));
        tmp(3385) := std_logic_vector(to_signed(-29062,16));
        tmp(3386) := std_logic_vector(to_signed(-29039,16));
        tmp(3387) := std_logic_vector(to_signed(-29016,16));
        tmp(3388) := std_logic_vector(to_signed(-28992,16));
        tmp(3389) := std_logic_vector(to_signed(-28969,16));
        tmp(3390) := std_logic_vector(to_signed(-28945,16));
        tmp(3391) := std_logic_vector(to_signed(-28922,16));
        tmp(3392) := std_logic_vector(to_signed(-28898,16));
        tmp(3393) := std_logic_vector(to_signed(-28874,16));
        tmp(3394) := std_logic_vector(to_signed(-28850,16));
        tmp(3395) := std_logic_vector(to_signed(-28827,16));
        tmp(3396) := std_logic_vector(to_signed(-28803,16));
        tmp(3397) := std_logic_vector(to_signed(-28779,16));
        tmp(3398) := std_logic_vector(to_signed(-28755,16));
        tmp(3399) := std_logic_vector(to_signed(-28730,16));
        tmp(3400) := std_logic_vector(to_signed(-28706,16));
        tmp(3401) := std_logic_vector(to_signed(-28682,16));
        tmp(3402) := std_logic_vector(to_signed(-28658,16));
        tmp(3403) := std_logic_vector(to_signed(-28633,16));
        tmp(3404) := std_logic_vector(to_signed(-28609,16));
        tmp(3405) := std_logic_vector(to_signed(-28584,16));
        tmp(3406) := std_logic_vector(to_signed(-28560,16));
        tmp(3407) := std_logic_vector(to_signed(-28535,16));
        tmp(3408) := std_logic_vector(to_signed(-28510,16));
        tmp(3409) := std_logic_vector(to_signed(-28485,16));
        tmp(3410) := std_logic_vector(to_signed(-28460,16));
        tmp(3411) := std_logic_vector(to_signed(-28436,16));
        tmp(3412) := std_logic_vector(to_signed(-28411,16));
        tmp(3413) := std_logic_vector(to_signed(-28385,16));
        tmp(3414) := std_logic_vector(to_signed(-28360,16));
        tmp(3415) := std_logic_vector(to_signed(-28335,16));
        tmp(3416) := std_logic_vector(to_signed(-28310,16));
        tmp(3417) := std_logic_vector(to_signed(-28284,16));
        tmp(3418) := std_logic_vector(to_signed(-28259,16));
        tmp(3419) := std_logic_vector(to_signed(-28234,16));
        tmp(3420) := std_logic_vector(to_signed(-28208,16));
        tmp(3421) := std_logic_vector(to_signed(-28182,16));
        tmp(3422) := std_logic_vector(to_signed(-28157,16));
        tmp(3423) := std_logic_vector(to_signed(-28131,16));
        tmp(3424) := std_logic_vector(to_signed(-28105,16));
        tmp(3425) := std_logic_vector(to_signed(-28079,16));
        tmp(3426) := std_logic_vector(to_signed(-28053,16));
        tmp(3427) := std_logic_vector(to_signed(-28027,16));
        tmp(3428) := std_logic_vector(to_signed(-28001,16));
        tmp(3429) := std_logic_vector(to_signed(-27975,16));
        tmp(3430) := std_logic_vector(to_signed(-27949,16));
        tmp(3431) := std_logic_vector(to_signed(-27923,16));
        tmp(3432) := std_logic_vector(to_signed(-27896,16));
        tmp(3433) := std_logic_vector(to_signed(-27870,16));
        tmp(3434) := std_logic_vector(to_signed(-27843,16));
        tmp(3435) := std_logic_vector(to_signed(-27817,16));
        tmp(3436) := std_logic_vector(to_signed(-27790,16));
        tmp(3437) := std_logic_vector(to_signed(-27764,16));
        tmp(3438) := std_logic_vector(to_signed(-27737,16));
        tmp(3439) := std_logic_vector(to_signed(-27710,16));
        tmp(3440) := std_logic_vector(to_signed(-27683,16));
        tmp(3441) := std_logic_vector(to_signed(-27656,16));
        tmp(3442) := std_logic_vector(to_signed(-27629,16));
        tmp(3443) := std_logic_vector(to_signed(-27602,16));
        tmp(3444) := std_logic_vector(to_signed(-27575,16));
        tmp(3445) := std_logic_vector(to_signed(-27548,16));
        tmp(3446) := std_logic_vector(to_signed(-27521,16));
        tmp(3447) := std_logic_vector(to_signed(-27493,16));
        tmp(3448) := std_logic_vector(to_signed(-27466,16));
        tmp(3449) := std_logic_vector(to_signed(-27439,16));
        tmp(3450) := std_logic_vector(to_signed(-27411,16));
        tmp(3451) := std_logic_vector(to_signed(-27384,16));
        tmp(3452) := std_logic_vector(to_signed(-27356,16));
        tmp(3453) := std_logic_vector(to_signed(-27328,16));
        tmp(3454) := std_logic_vector(to_signed(-27300,16));
        tmp(3455) := std_logic_vector(to_signed(-27273,16));
        tmp(3456) := std_logic_vector(to_signed(-27245,16));
        tmp(3457) := std_logic_vector(to_signed(-27217,16));
        tmp(3458) := std_logic_vector(to_signed(-27189,16));
        tmp(3459) := std_logic_vector(to_signed(-27161,16));
        tmp(3460) := std_logic_vector(to_signed(-27133,16));
        tmp(3461) := std_logic_vector(to_signed(-27104,16));
        tmp(3462) := std_logic_vector(to_signed(-27076,16));
        tmp(3463) := std_logic_vector(to_signed(-27048,16));
        tmp(3464) := std_logic_vector(to_signed(-27019,16));
        tmp(3465) := std_logic_vector(to_signed(-26991,16));
        tmp(3466) := std_logic_vector(to_signed(-26962,16));
        tmp(3467) := std_logic_vector(to_signed(-26934,16));
        tmp(3468) := std_logic_vector(to_signed(-26905,16));
        tmp(3469) := std_logic_vector(to_signed(-26876,16));
        tmp(3470) := std_logic_vector(to_signed(-26848,16));
        tmp(3471) := std_logic_vector(to_signed(-26819,16));
        tmp(3472) := std_logic_vector(to_signed(-26790,16));
        tmp(3473) := std_logic_vector(to_signed(-26761,16));
        tmp(3474) := std_logic_vector(to_signed(-26732,16));
        tmp(3475) := std_logic_vector(to_signed(-26703,16));
        tmp(3476) := std_logic_vector(to_signed(-26674,16));
        tmp(3477) := std_logic_vector(to_signed(-26644,16));
        tmp(3478) := std_logic_vector(to_signed(-26615,16));
        tmp(3479) := std_logic_vector(to_signed(-26586,16));
        tmp(3480) := std_logic_vector(to_signed(-26556,16));
        tmp(3481) := std_logic_vector(to_signed(-26527,16));
        tmp(3482) := std_logic_vector(to_signed(-26497,16));
        tmp(3483) := std_logic_vector(to_signed(-26468,16));
        tmp(3484) := std_logic_vector(to_signed(-26438,16));
        tmp(3485) := std_logic_vector(to_signed(-26408,16));
        tmp(3486) := std_logic_vector(to_signed(-26378,16));
        tmp(3487) := std_logic_vector(to_signed(-26349,16));
        tmp(3488) := std_logic_vector(to_signed(-26319,16));
        tmp(3489) := std_logic_vector(to_signed(-26289,16));
        tmp(3490) := std_logic_vector(to_signed(-26259,16));
        tmp(3491) := std_logic_vector(to_signed(-26229,16));
        tmp(3492) := std_logic_vector(to_signed(-26198,16));
        tmp(3493) := std_logic_vector(to_signed(-26168,16));
        tmp(3494) := std_logic_vector(to_signed(-26138,16));
        tmp(3495) := std_logic_vector(to_signed(-26108,16));
        tmp(3496) := std_logic_vector(to_signed(-26077,16));
        tmp(3497) := std_logic_vector(to_signed(-26047,16));
        tmp(3498) := std_logic_vector(to_signed(-26016,16));
        tmp(3499) := std_logic_vector(to_signed(-25986,16));
        tmp(3500) := std_logic_vector(to_signed(-25955,16));
        tmp(3501) := std_logic_vector(to_signed(-25924,16));
        tmp(3502) := std_logic_vector(to_signed(-25893,16));
        tmp(3503) := std_logic_vector(to_signed(-25863,16));
        tmp(3504) := std_logic_vector(to_signed(-25832,16));
        tmp(3505) := std_logic_vector(to_signed(-25801,16));
        tmp(3506) := std_logic_vector(to_signed(-25770,16));
        tmp(3507) := std_logic_vector(to_signed(-25739,16));
        tmp(3508) := std_logic_vector(to_signed(-25708,16));
        tmp(3509) := std_logic_vector(to_signed(-25676,16));
        tmp(3510) := std_logic_vector(to_signed(-25645,16));
        tmp(3511) := std_logic_vector(to_signed(-25614,16));
        tmp(3512) := std_logic_vector(to_signed(-25582,16));
        tmp(3513) := std_logic_vector(to_signed(-25551,16));
        tmp(3514) := std_logic_vector(to_signed(-25519,16));
        tmp(3515) := std_logic_vector(to_signed(-25488,16));
        tmp(3516) := std_logic_vector(to_signed(-25456,16));
        tmp(3517) := std_logic_vector(to_signed(-25425,16));
        tmp(3518) := std_logic_vector(to_signed(-25393,16));
        tmp(3519) := std_logic_vector(to_signed(-25361,16));
        tmp(3520) := std_logic_vector(to_signed(-25329,16));
        tmp(3521) := std_logic_vector(to_signed(-25297,16));
        tmp(3522) := std_logic_vector(to_signed(-25265,16));
        tmp(3523) := std_logic_vector(to_signed(-25233,16));
        tmp(3524) := std_logic_vector(to_signed(-25201,16));
        tmp(3525) := std_logic_vector(to_signed(-25169,16));
        tmp(3526) := std_logic_vector(to_signed(-25137,16));
        tmp(3527) := std_logic_vector(to_signed(-25105,16));
        tmp(3528) := std_logic_vector(to_signed(-25072,16));
        tmp(3529) := std_logic_vector(to_signed(-25040,16));
        tmp(3530) := std_logic_vector(to_signed(-25007,16));
        tmp(3531) := std_logic_vector(to_signed(-24975,16));
        tmp(3532) := std_logic_vector(to_signed(-24942,16));
        tmp(3533) := std_logic_vector(to_signed(-24910,16));
        tmp(3534) := std_logic_vector(to_signed(-24877,16));
        tmp(3535) := std_logic_vector(to_signed(-24844,16));
        tmp(3536) := std_logic_vector(to_signed(-24811,16));
        tmp(3537) := std_logic_vector(to_signed(-24779,16));
        tmp(3538) := std_logic_vector(to_signed(-24746,16));
        tmp(3539) := std_logic_vector(to_signed(-24713,16));
        tmp(3540) := std_logic_vector(to_signed(-24680,16));
        tmp(3541) := std_logic_vector(to_signed(-24647,16));
        tmp(3542) := std_logic_vector(to_signed(-24613,16));
        tmp(3543) := std_logic_vector(to_signed(-24580,16));
        tmp(3544) := std_logic_vector(to_signed(-24547,16));
        tmp(3545) := std_logic_vector(to_signed(-24514,16));
        tmp(3546) := std_logic_vector(to_signed(-24480,16));
        tmp(3547) := std_logic_vector(to_signed(-24447,16));
        tmp(3548) := std_logic_vector(to_signed(-24413,16));
        tmp(3549) := std_logic_vector(to_signed(-24380,16));
        tmp(3550) := std_logic_vector(to_signed(-24346,16));
        tmp(3551) := std_logic_vector(to_signed(-24312,16));
        tmp(3552) := std_logic_vector(to_signed(-24279,16));
        tmp(3553) := std_logic_vector(to_signed(-24245,16));
        tmp(3554) := std_logic_vector(to_signed(-24211,16));
        tmp(3555) := std_logic_vector(to_signed(-24177,16));
        tmp(3556) := std_logic_vector(to_signed(-24143,16));
        tmp(3557) := std_logic_vector(to_signed(-24109,16));
        tmp(3558) := std_logic_vector(to_signed(-24075,16));
        tmp(3559) := std_logic_vector(to_signed(-24041,16));
        tmp(3560) := std_logic_vector(to_signed(-24007,16));
        tmp(3561) := std_logic_vector(to_signed(-23973,16));
        tmp(3562) := std_logic_vector(to_signed(-23938,16));
        tmp(3563) := std_logic_vector(to_signed(-23904,16));
        tmp(3564) := std_logic_vector(to_signed(-23870,16));
        tmp(3565) := std_logic_vector(to_signed(-23835,16));
        tmp(3566) := std_logic_vector(to_signed(-23801,16));
        tmp(3567) := std_logic_vector(to_signed(-23766,16));
        tmp(3568) := std_logic_vector(to_signed(-23731,16));
        tmp(3569) := std_logic_vector(to_signed(-23697,16));
        tmp(3570) := std_logic_vector(to_signed(-23662,16));
        tmp(3571) := std_logic_vector(to_signed(-23627,16));
        tmp(3572) := std_logic_vector(to_signed(-23592,16));
        tmp(3573) := std_logic_vector(to_signed(-23557,16));
        tmp(3574) := std_logic_vector(to_signed(-23522,16));
        tmp(3575) := std_logic_vector(to_signed(-23487,16));
        tmp(3576) := std_logic_vector(to_signed(-23452,16));
        tmp(3577) := std_logic_vector(to_signed(-23417,16));
        tmp(3578) := std_logic_vector(to_signed(-23382,16));
        tmp(3579) := std_logic_vector(to_signed(-23347,16));
        tmp(3580) := std_logic_vector(to_signed(-23311,16));
        tmp(3581) := std_logic_vector(to_signed(-23276,16));
        tmp(3582) := std_logic_vector(to_signed(-23241,16));
        tmp(3583) := std_logic_vector(to_signed(-23205,16));
        tmp(3584) := std_logic_vector(to_signed(-23170,16));
        tmp(3585) := std_logic_vector(to_signed(-23134,16));
        tmp(3586) := std_logic_vector(to_signed(-23099,16));
        tmp(3587) := std_logic_vector(to_signed(-23063,16));
        tmp(3588) := std_logic_vector(to_signed(-23027,16));
        tmp(3589) := std_logic_vector(to_signed(-22991,16));
        tmp(3590) := std_logic_vector(to_signed(-22956,16));
        tmp(3591) := std_logic_vector(to_signed(-22920,16));
        tmp(3592) := std_logic_vector(to_signed(-22884,16));
        tmp(3593) := std_logic_vector(to_signed(-22848,16));
        tmp(3594) := std_logic_vector(to_signed(-22812,16));
        tmp(3595) := std_logic_vector(to_signed(-22776,16));
        tmp(3596) := std_logic_vector(to_signed(-22739,16));
        tmp(3597) := std_logic_vector(to_signed(-22703,16));
        tmp(3598) := std_logic_vector(to_signed(-22667,16));
        tmp(3599) := std_logic_vector(to_signed(-22631,16));
        tmp(3600) := std_logic_vector(to_signed(-22594,16));
        tmp(3601) := std_logic_vector(to_signed(-22558,16));
        tmp(3602) := std_logic_vector(to_signed(-22521,16));
        tmp(3603) := std_logic_vector(to_signed(-22485,16));
        tmp(3604) := std_logic_vector(to_signed(-22448,16));
        tmp(3605) := std_logic_vector(to_signed(-22411,16));
        tmp(3606) := std_logic_vector(to_signed(-22375,16));
        tmp(3607) := std_logic_vector(to_signed(-22338,16));
        tmp(3608) := std_logic_vector(to_signed(-22301,16));
        tmp(3609) := std_logic_vector(to_signed(-22264,16));
        tmp(3610) := std_logic_vector(to_signed(-22227,16));
        tmp(3611) := std_logic_vector(to_signed(-22191,16));
        tmp(3612) := std_logic_vector(to_signed(-22154,16));
        tmp(3613) := std_logic_vector(to_signed(-22116,16));
        tmp(3614) := std_logic_vector(to_signed(-22079,16));
        tmp(3615) := std_logic_vector(to_signed(-22042,16));
        tmp(3616) := std_logic_vector(to_signed(-22005,16));
        tmp(3617) := std_logic_vector(to_signed(-21968,16));
        tmp(3618) := std_logic_vector(to_signed(-21930,16));
        tmp(3619) := std_logic_vector(to_signed(-21893,16));
        tmp(3620) := std_logic_vector(to_signed(-21856,16));
        tmp(3621) := std_logic_vector(to_signed(-21818,16));
        tmp(3622) := std_logic_vector(to_signed(-21781,16));
        tmp(3623) := std_logic_vector(to_signed(-21743,16));
        tmp(3624) := std_logic_vector(to_signed(-21705,16));
        tmp(3625) := std_logic_vector(to_signed(-21668,16));
        tmp(3626) := std_logic_vector(to_signed(-21630,16));
        tmp(3627) := std_logic_vector(to_signed(-21592,16));
        tmp(3628) := std_logic_vector(to_signed(-21554,16));
        tmp(3629) := std_logic_vector(to_signed(-21516,16));
        tmp(3630) := std_logic_vector(to_signed(-21479,16));
        tmp(3631) := std_logic_vector(to_signed(-21441,16));
        tmp(3632) := std_logic_vector(to_signed(-21403,16));
        tmp(3633) := std_logic_vector(to_signed(-21364,16));
        tmp(3634) := std_logic_vector(to_signed(-21326,16));
        tmp(3635) := std_logic_vector(to_signed(-21288,16));
        tmp(3636) := std_logic_vector(to_signed(-21250,16));
        tmp(3637) := std_logic_vector(to_signed(-21212,16));
        tmp(3638) := std_logic_vector(to_signed(-21173,16));
        tmp(3639) := std_logic_vector(to_signed(-21135,16));
        tmp(3640) := std_logic_vector(to_signed(-21096,16));
        tmp(3641) := std_logic_vector(to_signed(-21058,16));
        tmp(3642) := std_logic_vector(to_signed(-21019,16));
        tmp(3643) := std_logic_vector(to_signed(-20981,16));
        tmp(3644) := std_logic_vector(to_signed(-20942,16));
        tmp(3645) := std_logic_vector(to_signed(-20904,16));
        tmp(3646) := std_logic_vector(to_signed(-20865,16));
        tmp(3647) := std_logic_vector(to_signed(-20826,16));
        tmp(3648) := std_logic_vector(to_signed(-20787,16));
        tmp(3649) := std_logic_vector(to_signed(-20748,16));
        tmp(3650) := std_logic_vector(to_signed(-20709,16));
        tmp(3651) := std_logic_vector(to_signed(-20670,16));
        tmp(3652) := std_logic_vector(to_signed(-20631,16));
        tmp(3653) := std_logic_vector(to_signed(-20592,16));
        tmp(3654) := std_logic_vector(to_signed(-20553,16));
        tmp(3655) := std_logic_vector(to_signed(-20514,16));
        tmp(3656) := std_logic_vector(to_signed(-20475,16));
        tmp(3657) := std_logic_vector(to_signed(-20436,16));
        tmp(3658) := std_logic_vector(to_signed(-20396,16));
        tmp(3659) := std_logic_vector(to_signed(-20357,16));
        tmp(3660) := std_logic_vector(to_signed(-20317,16));
        tmp(3661) := std_logic_vector(to_signed(-20278,16));
        tmp(3662) := std_logic_vector(to_signed(-20238,16));
        tmp(3663) := std_logic_vector(to_signed(-20199,16));
        tmp(3664) := std_logic_vector(to_signed(-20159,16));
        tmp(3665) := std_logic_vector(to_signed(-20120,16));
        tmp(3666) := std_logic_vector(to_signed(-20080,16));
        tmp(3667) := std_logic_vector(to_signed(-20040,16));
        tmp(3668) := std_logic_vector(to_signed(-20000,16));
        tmp(3669) := std_logic_vector(to_signed(-19961,16));
        tmp(3670) := std_logic_vector(to_signed(-19921,16));
        tmp(3671) := std_logic_vector(to_signed(-19881,16));
        tmp(3672) := std_logic_vector(to_signed(-19841,16));
        tmp(3673) := std_logic_vector(to_signed(-19801,16));
        tmp(3674) := std_logic_vector(to_signed(-19761,16));
        tmp(3675) := std_logic_vector(to_signed(-19721,16));
        tmp(3676) := std_logic_vector(to_signed(-19680,16));
        tmp(3677) := std_logic_vector(to_signed(-19640,16));
        tmp(3678) := std_logic_vector(to_signed(-19600,16));
        tmp(3679) := std_logic_vector(to_signed(-19560,16));
        tmp(3680) := std_logic_vector(to_signed(-19519,16));
        tmp(3681) := std_logic_vector(to_signed(-19479,16));
        tmp(3682) := std_logic_vector(to_signed(-19438,16));
        tmp(3683) := std_logic_vector(to_signed(-19398,16));
        tmp(3684) := std_logic_vector(to_signed(-19357,16));
        tmp(3685) := std_logic_vector(to_signed(-19317,16));
        tmp(3686) := std_logic_vector(to_signed(-19276,16));
        tmp(3687) := std_logic_vector(to_signed(-19236,16));
        tmp(3688) := std_logic_vector(to_signed(-19195,16));
        tmp(3689) := std_logic_vector(to_signed(-19154,16));
        tmp(3690) := std_logic_vector(to_signed(-19113,16));
        tmp(3691) := std_logic_vector(to_signed(-19072,16));
        tmp(3692) := std_logic_vector(to_signed(-19032,16));
        tmp(3693) := std_logic_vector(to_signed(-18991,16));
        tmp(3694) := std_logic_vector(to_signed(-18950,16));
        tmp(3695) := std_logic_vector(to_signed(-18909,16));
        tmp(3696) := std_logic_vector(to_signed(-18868,16));
        tmp(3697) := std_logic_vector(to_signed(-18826,16));
        tmp(3698) := std_logic_vector(to_signed(-18785,16));
        tmp(3699) := std_logic_vector(to_signed(-18744,16));
        tmp(3700) := std_logic_vector(to_signed(-18703,16));
        tmp(3701) := std_logic_vector(to_signed(-18661,16));
        tmp(3702) := std_logic_vector(to_signed(-18620,16));
        tmp(3703) := std_logic_vector(to_signed(-18579,16));
        tmp(3704) := std_logic_vector(to_signed(-18537,16));
        tmp(3705) := std_logic_vector(to_signed(-18496,16));
        tmp(3706) := std_logic_vector(to_signed(-18454,16));
        tmp(3707) := std_logic_vector(to_signed(-18413,16));
        tmp(3708) := std_logic_vector(to_signed(-18371,16));
        tmp(3709) := std_logic_vector(to_signed(-18330,16));
        tmp(3710) := std_logic_vector(to_signed(-18288,16));
        tmp(3711) := std_logic_vector(to_signed(-18246,16));
        tmp(3712) := std_logic_vector(to_signed(-18204,16));
        tmp(3713) := std_logic_vector(to_signed(-18163,16));
        tmp(3714) := std_logic_vector(to_signed(-18121,16));
        tmp(3715) := std_logic_vector(to_signed(-18079,16));
        tmp(3716) := std_logic_vector(to_signed(-18037,16));
        tmp(3717) := std_logic_vector(to_signed(-17995,16));
        tmp(3718) := std_logic_vector(to_signed(-17953,16));
        tmp(3719) := std_logic_vector(to_signed(-17911,16));
        tmp(3720) := std_logic_vector(to_signed(-17869,16));
        tmp(3721) := std_logic_vector(to_signed(-17827,16));
        tmp(3722) := std_logic_vector(to_signed(-17784,16));
        tmp(3723) := std_logic_vector(to_signed(-17742,16));
        tmp(3724) := std_logic_vector(to_signed(-17700,16));
        tmp(3725) := std_logic_vector(to_signed(-17657,16));
        tmp(3726) := std_logic_vector(to_signed(-17615,16));
        tmp(3727) := std_logic_vector(to_signed(-17573,16));
        tmp(3728) := std_logic_vector(to_signed(-17530,16));
        tmp(3729) := std_logic_vector(to_signed(-17488,16));
        tmp(3730) := std_logic_vector(to_signed(-17445,16));
        tmp(3731) := std_logic_vector(to_signed(-17403,16));
        tmp(3732) := std_logic_vector(to_signed(-17360,16));
        tmp(3733) := std_logic_vector(to_signed(-17317,16));
        tmp(3734) := std_logic_vector(to_signed(-17275,16));
        tmp(3735) := std_logic_vector(to_signed(-17232,16));
        tmp(3736) := std_logic_vector(to_signed(-17189,16));
        tmp(3737) := std_logic_vector(to_signed(-17146,16));
        tmp(3738) := std_logic_vector(to_signed(-17104,16));
        tmp(3739) := std_logic_vector(to_signed(-17061,16));
        tmp(3740) := std_logic_vector(to_signed(-17018,16));
        tmp(3741) := std_logic_vector(to_signed(-16975,16));
        tmp(3742) := std_logic_vector(to_signed(-16932,16));
        tmp(3743) := std_logic_vector(to_signed(-16889,16));
        tmp(3744) := std_logic_vector(to_signed(-16846,16));
        tmp(3745) := std_logic_vector(to_signed(-16802,16));
        tmp(3746) := std_logic_vector(to_signed(-16759,16));
        tmp(3747) := std_logic_vector(to_signed(-16716,16));
        tmp(3748) := std_logic_vector(to_signed(-16673,16));
        tmp(3749) := std_logic_vector(to_signed(-16630,16));
        tmp(3750) := std_logic_vector(to_signed(-16586,16));
        tmp(3751) := std_logic_vector(to_signed(-16543,16));
        tmp(3752) := std_logic_vector(to_signed(-16499,16));
        tmp(3753) := std_logic_vector(to_signed(-16456,16));
        tmp(3754) := std_logic_vector(to_signed(-16413,16));
        tmp(3755) := std_logic_vector(to_signed(-16369,16));
        tmp(3756) := std_logic_vector(to_signed(-16325,16));
        tmp(3757) := std_logic_vector(to_signed(-16282,16));
        tmp(3758) := std_logic_vector(to_signed(-16238,16));
        tmp(3759) := std_logic_vector(to_signed(-16195,16));
        tmp(3760) := std_logic_vector(to_signed(-16151,16));
        tmp(3761) := std_logic_vector(to_signed(-16107,16));
        tmp(3762) := std_logic_vector(to_signed(-16063,16));
        tmp(3763) := std_logic_vector(to_signed(-16019,16));
        tmp(3764) := std_logic_vector(to_signed(-15976,16));
        tmp(3765) := std_logic_vector(to_signed(-15932,16));
        tmp(3766) := std_logic_vector(to_signed(-15888,16));
        tmp(3767) := std_logic_vector(to_signed(-15844,16));
        tmp(3768) := std_logic_vector(to_signed(-15800,16));
        tmp(3769) := std_logic_vector(to_signed(-15756,16));
        tmp(3770) := std_logic_vector(to_signed(-15712,16));
        tmp(3771) := std_logic_vector(to_signed(-15667,16));
        tmp(3772) := std_logic_vector(to_signed(-15623,16));
        tmp(3773) := std_logic_vector(to_signed(-15579,16));
        tmp(3774) := std_logic_vector(to_signed(-15535,16));
        tmp(3775) := std_logic_vector(to_signed(-15491,16));
        tmp(3776) := std_logic_vector(to_signed(-15446,16));
        tmp(3777) := std_logic_vector(to_signed(-15402,16));
        tmp(3778) := std_logic_vector(to_signed(-15358,16));
        tmp(3779) := std_logic_vector(to_signed(-15313,16));
        tmp(3780) := std_logic_vector(to_signed(-15269,16));
        tmp(3781) := std_logic_vector(to_signed(-15224,16));
        tmp(3782) := std_logic_vector(to_signed(-15180,16));
        tmp(3783) := std_logic_vector(to_signed(-15135,16));
        tmp(3784) := std_logic_vector(to_signed(-15090,16));
        tmp(3785) := std_logic_vector(to_signed(-15046,16));
        tmp(3786) := std_logic_vector(to_signed(-15001,16));
        tmp(3787) := std_logic_vector(to_signed(-14956,16));
        tmp(3788) := std_logic_vector(to_signed(-14912,16));
        tmp(3789) := std_logic_vector(to_signed(-14867,16));
        tmp(3790) := std_logic_vector(to_signed(-14822,16));
        tmp(3791) := std_logic_vector(to_signed(-14777,16));
        tmp(3792) := std_logic_vector(to_signed(-14732,16));
        tmp(3793) := std_logic_vector(to_signed(-14688,16));
        tmp(3794) := std_logic_vector(to_signed(-14643,16));
        tmp(3795) := std_logic_vector(to_signed(-14598,16));
        tmp(3796) := std_logic_vector(to_signed(-14553,16));
        tmp(3797) := std_logic_vector(to_signed(-14507,16));
        tmp(3798) := std_logic_vector(to_signed(-14462,16));
        tmp(3799) := std_logic_vector(to_signed(-14417,16));
        tmp(3800) := std_logic_vector(to_signed(-14372,16));
        tmp(3801) := std_logic_vector(to_signed(-14327,16));
        tmp(3802) := std_logic_vector(to_signed(-14282,16));
        tmp(3803) := std_logic_vector(to_signed(-14236,16));
        tmp(3804) := std_logic_vector(to_signed(-14191,16));
        tmp(3805) := std_logic_vector(to_signed(-14146,16));
        tmp(3806) := std_logic_vector(to_signed(-14101,16));
        tmp(3807) := std_logic_vector(to_signed(-14055,16));
        tmp(3808) := std_logic_vector(to_signed(-14010,16));
        tmp(3809) := std_logic_vector(to_signed(-13964,16));
        tmp(3810) := std_logic_vector(to_signed(-13919,16));
        tmp(3811) := std_logic_vector(to_signed(-13873,16));
        tmp(3812) := std_logic_vector(to_signed(-13828,16));
        tmp(3813) := std_logic_vector(to_signed(-13782,16));
        tmp(3814) := std_logic_vector(to_signed(-13736,16));
        tmp(3815) := std_logic_vector(to_signed(-13691,16));
        tmp(3816) := std_logic_vector(to_signed(-13645,16));
        tmp(3817) := std_logic_vector(to_signed(-13599,16));
        tmp(3818) := std_logic_vector(to_signed(-13554,16));
        tmp(3819) := std_logic_vector(to_signed(-13508,16));
        tmp(3820) := std_logic_vector(to_signed(-13462,16));
        tmp(3821) := std_logic_vector(to_signed(-13416,16));
        tmp(3822) := std_logic_vector(to_signed(-13370,16));
        tmp(3823) := std_logic_vector(to_signed(-13324,16));
        tmp(3824) := std_logic_vector(to_signed(-13279,16));
        tmp(3825) := std_logic_vector(to_signed(-13233,16));
        tmp(3826) := std_logic_vector(to_signed(-13187,16));
        tmp(3827) := std_logic_vector(to_signed(-13141,16));
        tmp(3828) := std_logic_vector(to_signed(-13094,16));
        tmp(3829) := std_logic_vector(to_signed(-13048,16));
        tmp(3830) := std_logic_vector(to_signed(-13002,16));
        tmp(3831) := std_logic_vector(to_signed(-12956,16));
        tmp(3832) := std_logic_vector(to_signed(-12910,16));
        tmp(3833) := std_logic_vector(to_signed(-12864,16));
        tmp(3834) := std_logic_vector(to_signed(-12817,16));
        tmp(3835) := std_logic_vector(to_signed(-12771,16));
        tmp(3836) := std_logic_vector(to_signed(-12725,16));
        tmp(3837) := std_logic_vector(to_signed(-12679,16));
        tmp(3838) := std_logic_vector(to_signed(-12632,16));
        tmp(3839) := std_logic_vector(to_signed(-12586,16));
        tmp(3840) := std_logic_vector(to_signed(-12539,16));
        tmp(3841) := std_logic_vector(to_signed(-12493,16));
        tmp(3842) := std_logic_vector(to_signed(-12446,16));
        tmp(3843) := std_logic_vector(to_signed(-12400,16));
        tmp(3844) := std_logic_vector(to_signed(-12353,16));
        tmp(3845) := std_logic_vector(to_signed(-12307,16));
        tmp(3846) := std_logic_vector(to_signed(-12260,16));
        tmp(3847) := std_logic_vector(to_signed(-12214,16));
        tmp(3848) := std_logic_vector(to_signed(-12167,16));
        tmp(3849) := std_logic_vector(to_signed(-12120,16));
        tmp(3850) := std_logic_vector(to_signed(-12074,16));
        tmp(3851) := std_logic_vector(to_signed(-12027,16));
        tmp(3852) := std_logic_vector(to_signed(-11980,16));
        tmp(3853) := std_logic_vector(to_signed(-11933,16));
        tmp(3854) := std_logic_vector(to_signed(-11886,16));
        tmp(3855) := std_logic_vector(to_signed(-11840,16));
        tmp(3856) := std_logic_vector(to_signed(-11793,16));
        tmp(3857) := std_logic_vector(to_signed(-11746,16));
        tmp(3858) := std_logic_vector(to_signed(-11699,16));
        tmp(3859) := std_logic_vector(to_signed(-11652,16));
        tmp(3860) := std_logic_vector(to_signed(-11605,16));
        tmp(3861) := std_logic_vector(to_signed(-11558,16));
        tmp(3862) := std_logic_vector(to_signed(-11511,16));
        tmp(3863) := std_logic_vector(to_signed(-11464,16));
        tmp(3864) := std_logic_vector(to_signed(-11417,16));
        tmp(3865) := std_logic_vector(to_signed(-11370,16));
        tmp(3866) := std_logic_vector(to_signed(-11322,16));
        tmp(3867) := std_logic_vector(to_signed(-11275,16));
        tmp(3868) := std_logic_vector(to_signed(-11228,16));
        tmp(3869) := std_logic_vector(to_signed(-11181,16));
        tmp(3870) := std_logic_vector(to_signed(-11133,16));
        tmp(3871) := std_logic_vector(to_signed(-11086,16));
        tmp(3872) := std_logic_vector(to_signed(-11039,16));
        tmp(3873) := std_logic_vector(to_signed(-10992,16));
        tmp(3874) := std_logic_vector(to_signed(-10944,16));
        tmp(3875) := std_logic_vector(to_signed(-10897,16));
        tmp(3876) := std_logic_vector(to_signed(-10849,16));
        tmp(3877) := std_logic_vector(to_signed(-10802,16));
        tmp(3878) := std_logic_vector(to_signed(-10754,16));
        tmp(3879) := std_logic_vector(to_signed(-10707,16));
        tmp(3880) := std_logic_vector(to_signed(-10659,16));
        tmp(3881) := std_logic_vector(to_signed(-10612,16));
        tmp(3882) := std_logic_vector(to_signed(-10564,16));
        tmp(3883) := std_logic_vector(to_signed(-10517,16));
        tmp(3884) := std_logic_vector(to_signed(-10469,16));
        tmp(3885) := std_logic_vector(to_signed(-10421,16));
        tmp(3886) := std_logic_vector(to_signed(-10374,16));
        tmp(3887) := std_logic_vector(to_signed(-10326,16));
        tmp(3888) := std_logic_vector(to_signed(-10278,16));
        tmp(3889) := std_logic_vector(to_signed(-10231,16));
        tmp(3890) := std_logic_vector(to_signed(-10183,16));
        tmp(3891) := std_logic_vector(to_signed(-10135,16));
        tmp(3892) := std_logic_vector(to_signed(-10087,16));
        tmp(3893) := std_logic_vector(to_signed(-10039,16));
        tmp(3894) := std_logic_vector(to_signed(-9992,16));
        tmp(3895) := std_logic_vector(to_signed(-9944,16));
        tmp(3896) := std_logic_vector(to_signed(-9896,16));
        tmp(3897) := std_logic_vector(to_signed(-9848,16));
        tmp(3898) := std_logic_vector(to_signed(-9800,16));
        tmp(3899) := std_logic_vector(to_signed(-9752,16));
        tmp(3900) := std_logic_vector(to_signed(-9704,16));
        tmp(3901) := std_logic_vector(to_signed(-9656,16));
        tmp(3902) := std_logic_vector(to_signed(-9608,16));
        tmp(3903) := std_logic_vector(to_signed(-9560,16));
        tmp(3904) := std_logic_vector(to_signed(-9512,16));
        tmp(3905) := std_logic_vector(to_signed(-9464,16));
        tmp(3906) := std_logic_vector(to_signed(-9416,16));
        tmp(3907) := std_logic_vector(to_signed(-9367,16));
        tmp(3908) := std_logic_vector(to_signed(-9319,16));
        tmp(3909) := std_logic_vector(to_signed(-9271,16));
        tmp(3910) := std_logic_vector(to_signed(-9223,16));
        tmp(3911) := std_logic_vector(to_signed(-9175,16));
        tmp(3912) := std_logic_vector(to_signed(-9126,16));
        tmp(3913) := std_logic_vector(to_signed(-9078,16));
        tmp(3914) := std_logic_vector(to_signed(-9030,16));
        tmp(3915) := std_logic_vector(to_signed(-8981,16));
        tmp(3916) := std_logic_vector(to_signed(-8933,16));
        tmp(3917) := std_logic_vector(to_signed(-8885,16));
        tmp(3918) := std_logic_vector(to_signed(-8836,16));
        tmp(3919) := std_logic_vector(to_signed(-8788,16));
        tmp(3920) := std_logic_vector(to_signed(-8739,16));
        tmp(3921) := std_logic_vector(to_signed(-8691,16));
        tmp(3922) := std_logic_vector(to_signed(-8642,16));
        tmp(3923) := std_logic_vector(to_signed(-8594,16));
        tmp(3924) := std_logic_vector(to_signed(-8545,16));
        tmp(3925) := std_logic_vector(to_signed(-8497,16));
        tmp(3926) := std_logic_vector(to_signed(-8448,16));
        tmp(3927) := std_logic_vector(to_signed(-8400,16));
        tmp(3928) := std_logic_vector(to_signed(-8351,16));
        tmp(3929) := std_logic_vector(to_signed(-8303,16));
        tmp(3930) := std_logic_vector(to_signed(-8254,16));
        tmp(3931) := std_logic_vector(to_signed(-8205,16));
        tmp(3932) := std_logic_vector(to_signed(-8157,16));
        tmp(3933) := std_logic_vector(to_signed(-8108,16));
        tmp(3934) := std_logic_vector(to_signed(-8059,16));
        tmp(3935) := std_logic_vector(to_signed(-8010,16));
        tmp(3936) := std_logic_vector(to_signed(-7962,16));
        tmp(3937) := std_logic_vector(to_signed(-7913,16));
        tmp(3938) := std_logic_vector(to_signed(-7864,16));
        tmp(3939) := std_logic_vector(to_signed(-7815,16));
        tmp(3940) := std_logic_vector(to_signed(-7767,16));
        tmp(3941) := std_logic_vector(to_signed(-7718,16));
        tmp(3942) := std_logic_vector(to_signed(-7669,16));
        tmp(3943) := std_logic_vector(to_signed(-7620,16));
        tmp(3944) := std_logic_vector(to_signed(-7571,16));
        tmp(3945) := std_logic_vector(to_signed(-7522,16));
        tmp(3946) := std_logic_vector(to_signed(-7473,16));
        tmp(3947) := std_logic_vector(to_signed(-7424,16));
        tmp(3948) := std_logic_vector(to_signed(-7375,16));
        tmp(3949) := std_logic_vector(to_signed(-7326,16));
        tmp(3950) := std_logic_vector(to_signed(-7277,16));
        tmp(3951) := std_logic_vector(to_signed(-7228,16));
        tmp(3952) := std_logic_vector(to_signed(-7179,16));
        tmp(3953) := std_logic_vector(to_signed(-7130,16));
        tmp(3954) := std_logic_vector(to_signed(-7081,16));
        tmp(3955) := std_logic_vector(to_signed(-7032,16));
        tmp(3956) := std_logic_vector(to_signed(-6983,16));
        tmp(3957) := std_logic_vector(to_signed(-6934,16));
        tmp(3958) := std_logic_vector(to_signed(-6885,16));
        tmp(3959) := std_logic_vector(to_signed(-6836,16));
        tmp(3960) := std_logic_vector(to_signed(-6786,16));
        tmp(3961) := std_logic_vector(to_signed(-6737,16));
        tmp(3962) := std_logic_vector(to_signed(-6688,16));
        tmp(3963) := std_logic_vector(to_signed(-6639,16));
        tmp(3964) := std_logic_vector(to_signed(-6590,16));
        tmp(3965) := std_logic_vector(to_signed(-6540,16));
        tmp(3966) := std_logic_vector(to_signed(-6491,16));
        tmp(3967) := std_logic_vector(to_signed(-6442,16));
        tmp(3968) := std_logic_vector(to_signed(-6393,16));
        tmp(3969) := std_logic_vector(to_signed(-6343,16));
        tmp(3970) := std_logic_vector(to_signed(-6294,16));
        tmp(3971) := std_logic_vector(to_signed(-6245,16));
        tmp(3972) := std_logic_vector(to_signed(-6195,16));
        tmp(3973) := std_logic_vector(to_signed(-6146,16));
        tmp(3974) := std_logic_vector(to_signed(-6096,16));
        tmp(3975) := std_logic_vector(to_signed(-6047,16));
        tmp(3976) := std_logic_vector(to_signed(-5998,16));
        tmp(3977) := std_logic_vector(to_signed(-5948,16));
        tmp(3978) := std_logic_vector(to_signed(-5899,16));
        tmp(3979) := std_logic_vector(to_signed(-5849,16));
        tmp(3980) := std_logic_vector(to_signed(-5800,16));
        tmp(3981) := std_logic_vector(to_signed(-5750,16));
        tmp(3982) := std_logic_vector(to_signed(-5701,16));
        tmp(3983) := std_logic_vector(to_signed(-5651,16));
        tmp(3984) := std_logic_vector(to_signed(-5602,16));
        tmp(3985) := std_logic_vector(to_signed(-5552,16));
        tmp(3986) := std_logic_vector(to_signed(-5503,16));
        tmp(3987) := std_logic_vector(to_signed(-5453,16));
        tmp(3988) := std_logic_vector(to_signed(-5404,16));
        tmp(3989) := std_logic_vector(to_signed(-5354,16));
        tmp(3990) := std_logic_vector(to_signed(-5305,16));
        tmp(3991) := std_logic_vector(to_signed(-5255,16));
        tmp(3992) := std_logic_vector(to_signed(-5205,16));
        tmp(3993) := std_logic_vector(to_signed(-5156,16));
        tmp(3994) := std_logic_vector(to_signed(-5106,16));
        tmp(3995) := std_logic_vector(to_signed(-5056,16));
        tmp(3996) := std_logic_vector(to_signed(-5007,16));
        tmp(3997) := std_logic_vector(to_signed(-4957,16));
        tmp(3998) := std_logic_vector(to_signed(-4907,16));
        tmp(3999) := std_logic_vector(to_signed(-4858,16));
        tmp(4000) := std_logic_vector(to_signed(-4808,16));
        tmp(4001) := std_logic_vector(to_signed(-4758,16));
        tmp(4002) := std_logic_vector(to_signed(-4708,16));
        tmp(4003) := std_logic_vector(to_signed(-4659,16));
        tmp(4004) := std_logic_vector(to_signed(-4609,16));
        tmp(4005) := std_logic_vector(to_signed(-4559,16));
        tmp(4006) := std_logic_vector(to_signed(-4509,16));
        tmp(4007) := std_logic_vector(to_signed(-4460,16));
        tmp(4008) := std_logic_vector(to_signed(-4410,16));
        tmp(4009) := std_logic_vector(to_signed(-4360,16));
        tmp(4010) := std_logic_vector(to_signed(-4310,16));
        tmp(4011) := std_logic_vector(to_signed(-4260,16));
        tmp(4012) := std_logic_vector(to_signed(-4210,16));
        tmp(4013) := std_logic_vector(to_signed(-4161,16));
        tmp(4014) := std_logic_vector(to_signed(-4111,16));
        tmp(4015) := std_logic_vector(to_signed(-4061,16));
        tmp(4016) := std_logic_vector(to_signed(-4011,16));
        tmp(4017) := std_logic_vector(to_signed(-3961,16));
        tmp(4018) := std_logic_vector(to_signed(-3911,16));
        tmp(4019) := std_logic_vector(to_signed(-3861,16));
        tmp(4020) := std_logic_vector(to_signed(-3811,16));
        tmp(4021) := std_logic_vector(to_signed(-3761,16));
        tmp(4022) := std_logic_vector(to_signed(-3712,16));
        tmp(4023) := std_logic_vector(to_signed(-3662,16));
        tmp(4024) := std_logic_vector(to_signed(-3612,16));
        tmp(4025) := std_logic_vector(to_signed(-3562,16));
        tmp(4026) := std_logic_vector(to_signed(-3512,16));
        tmp(4027) := std_logic_vector(to_signed(-3462,16));
        tmp(4028) := std_logic_vector(to_signed(-3412,16));
        tmp(4029) := std_logic_vector(to_signed(-3362,16));
        tmp(4030) := std_logic_vector(to_signed(-3312,16));
        tmp(4031) := std_logic_vector(to_signed(-3262,16));
        tmp(4032) := std_logic_vector(to_signed(-3212,16));
        tmp(4033) := std_logic_vector(to_signed(-3162,16));
        tmp(4034) := std_logic_vector(to_signed(-3112,16));
        tmp(4035) := std_logic_vector(to_signed(-3062,16));
        tmp(4036) := std_logic_vector(to_signed(-3012,16));
        tmp(4037) := std_logic_vector(to_signed(-2962,16));
        tmp(4038) := std_logic_vector(to_signed(-2911,16));
        tmp(4039) := std_logic_vector(to_signed(-2861,16));
        tmp(4040) := std_logic_vector(to_signed(-2811,16));
        tmp(4041) := std_logic_vector(to_signed(-2761,16));
        tmp(4042) := std_logic_vector(to_signed(-2711,16));
        tmp(4043) := std_logic_vector(to_signed(-2661,16));
        tmp(4044) := std_logic_vector(to_signed(-2611,16));
        tmp(4045) := std_logic_vector(to_signed(-2561,16));
        tmp(4046) := std_logic_vector(to_signed(-2511,16));
        tmp(4047) := std_logic_vector(to_signed(-2461,16));
        tmp(4048) := std_logic_vector(to_signed(-2410,16));
        tmp(4049) := std_logic_vector(to_signed(-2360,16));
        tmp(4050) := std_logic_vector(to_signed(-2310,16));
        tmp(4051) := std_logic_vector(to_signed(-2260,16));
        tmp(4052) := std_logic_vector(to_signed(-2210,16));
        tmp(4053) := std_logic_vector(to_signed(-2160,16));
        tmp(4054) := std_logic_vector(to_signed(-2110,16));
        tmp(4055) := std_logic_vector(to_signed(-2059,16));
        tmp(4056) := std_logic_vector(to_signed(-2009,16));
        tmp(4057) := std_logic_vector(to_signed(-1959,16));
        tmp(4058) := std_logic_vector(to_signed(-1909,16));
        tmp(4059) := std_logic_vector(to_signed(-1859,16));
        tmp(4060) := std_logic_vector(to_signed(-1809,16));
        tmp(4061) := std_logic_vector(to_signed(-1758,16));
        tmp(4062) := std_logic_vector(to_signed(-1708,16));
        tmp(4063) := std_logic_vector(to_signed(-1658,16));
        tmp(4064) := std_logic_vector(to_signed(-1608,16));
        tmp(4065) := std_logic_vector(to_signed(-1558,16));
        tmp(4066) := std_logic_vector(to_signed(-1507,16));
        tmp(4067) := std_logic_vector(to_signed(-1457,16));
        tmp(4068) := std_logic_vector(to_signed(-1407,16));
        tmp(4069) := std_logic_vector(to_signed(-1357,16));
        tmp(4070) := std_logic_vector(to_signed(-1307,16));
        tmp(4071) := std_logic_vector(to_signed(-1256,16));
        tmp(4072) := std_logic_vector(to_signed(-1206,16));
        tmp(4073) := std_logic_vector(to_signed(-1156,16));
        tmp(4074) := std_logic_vector(to_signed(-1106,16));
        tmp(4075) := std_logic_vector(to_signed(-1055,16));
        tmp(4076) := std_logic_vector(to_signed(-1005,16));
        tmp(4077) := std_logic_vector(to_signed(-955,16));
        tmp(4078) := std_logic_vector(to_signed(-905,16));
        tmp(4079) := std_logic_vector(to_signed(-854,16));
        tmp(4080) := std_logic_vector(to_signed(-804,16));
        tmp(4081) := std_logic_vector(to_signed(-754,16));
        tmp(4082) := std_logic_vector(to_signed(-704,16));
        tmp(4083) := std_logic_vector(to_signed(-653,16));
        tmp(4084) := std_logic_vector(to_signed(-603,16));
        tmp(4085) := std_logic_vector(to_signed(-553,16));
        tmp(4086) := std_logic_vector(to_signed(-503,16));
        tmp(4087) := std_logic_vector(to_signed(-452,16));
        tmp(4088) := std_logic_vector(to_signed(-402,16));
        tmp(4089) := std_logic_vector(to_signed(-352,16));
        tmp(4090) := std_logic_vector(to_signed(-302,16));
        tmp(4091) := std_logic_vector(to_signed(-251,16));
        tmp(4092) := std_logic_vector(to_signed(-201,16));
        tmp(4093) := std_logic_vector(to_signed(-151,16));
        tmp(4094) := std_logic_vector(to_signed(-101,16));
        tmp(4095) := std_logic_vector(to_signed(-50,16));
	return tmp;                                                              
end init_rom;                                                               
signal ROM: ROM_type:=init_rom;                                                         
                                                                              
begin                                                                         
                                                                              
process(clk)                                                                  
begin                                                                         
    if rising_edge(clk) then                                                  
            data_out <= ROM(to_integer(unsigned(addr_in)));                                           
    end if;                                                                   
end process;                                                                  
                                                                              
end rtl;                                                                      
