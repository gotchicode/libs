library IEEE;                                                                                                                            
use IEEE.std_logic_1164.all;                                                                                                             
use IEEE.numeric_std.all;                                                                                                                
                                                                                                                                         
entity top is                                                                                                                            
 port (                                                                                                                                  
            clk             : in std_logic;                                                                                              
                                                                                                                                         
            data_in         : in std_logic;                                                                                              
			data_out		: out std_logic_vector(3 downto 0)                                                                            
                                                                                                                                         
 );                                                                                                                                      
end entity top;                                                                                                                          
                                                                                                                                         
architecture rtl of top is                                                                                                               
                                                                                                                                         
constant USE_MITIGATION             : integer:=0;                                                                                        
                                                                                                                                         
constant nb_reg                     : integer:=1000; --(nb_reg-1 LUT on Xilinx target without mitigation)                                  
                                                                                                                                         
--signal lut_in                   : std_logic_vector(nb_reg-1 downto 0);                                                                 
--signal lut_out                  : std_logic_vector(nb_reg-1 downto 0);                                                                 
                                                                                                                                         
signal registers                    : std_logic_vector(nb_reg-1 downto 0);                                                               
--signal registers_d1             : std_logic_vector(nb_reg-1 downto 0);                                                                 
                                                                                                                                         
type tmr_reg_type                   is array (0 to 2) of std_logic_vector(nb_reg-1 downto 0);                                            
signal tmr_registers                : tmr_reg_type;                                                                                      
signal local_tmr_voter              : std_logic_vector(nb_reg-1 downto 0);                                                               
signal global_tmr_voter             : tmr_reg_type;                                                                                      
                                                                                                                                         
attribute keep                      : string;                                                                                            
attribute keep of registers         : signal is "true";                                                                                  
attribute keep of tmr_registers     : signal is "true";                                                                                  
attribute keep of local_tmr_voter   : signal is "true";                                                                                  
attribute keep of global_tmr_voter  : signal is "true";                                                                                  
-- synthesis translate_on 
attribute syn_keep of registers, tmr_registers, local_tmr_voter, global_tmr_voter : signal is true;
-- synthesis translate_off 
                                                                                                                                         
begin                                                                                                                                    
                                                                                                                                         
----------------------------------------------------------------------------------------------------------------------------             
--                                                                                                                                       
--                                                                                                                                       
--              NO MITIGATION IN THE DESIGN                                                                                              
--                                                                                                                                       
--                                                                                                                                       
----------------------------------------------------------------------------------------------------------------------------             
                                                                                                                                         
NO_MITIGATION: if USE_MITIGATION=0 generate                                                                                              
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Input                                                                                                                             
    ------------------------------------------                                                                                           
    registers(0) <= data_in;                                                                                                             
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Combinatiorial + Registers                                                                                                        
    ------------------------------------------                                                                                           
    process(clk)                                                                                                                         
    begin                                                                                                                                
                                                                                                                                         
        if rising_edge(clk) then                                                                                                         
                                                                                                                                         
                registers(1)    <= not(registers(0));                                                                              
                registers(2)    <= not(registers(1));                                                                              
                registers(3)    <= not(registers(2));                                                                              
                registers(4)    <= not(registers(3));                                                                              
                registers(5)    <= not(registers(4));                                                                              
                registers(6)    <= not(registers(5));                                                                              
                registers(7)    <= not(registers(6));                                                                              
                registers(8)    <= not(registers(7));                                                                              
                registers(9)    <= not(registers(8));                                                                              
                registers(10)    <= not(registers(9));                                                                              
                registers(11)    <= not(registers(10));                                                                              
                registers(12)    <= not(registers(11));                                                                              
                registers(13)    <= not(registers(12));                                                                              
                registers(14)    <= not(registers(13));                                                                              
                registers(15)    <= not(registers(14));                                                                              
                registers(16)    <= not(registers(15));                                                                              
                registers(17)    <= not(registers(16));                                                                              
                registers(18)    <= not(registers(17));                                                                              
                registers(19)    <= not(registers(18));                                                                              
                registers(20)    <= not(registers(19));                                                                              
                registers(21)    <= not(registers(20));                                                                              
                registers(22)    <= not(registers(21));                                                                              
                registers(23)    <= not(registers(22));                                                                              
                registers(24)    <= not(registers(23));                                                                              
                registers(25)    <= not(registers(24));                                                                              
                registers(26)    <= not(registers(25));                                                                              
                registers(27)    <= not(registers(26));                                                                              
                registers(28)    <= not(registers(27));                                                                              
                registers(29)    <= not(registers(28));                                                                              
                registers(30)    <= not(registers(29));                                                                              
                registers(31)    <= not(registers(30));                                                                              
                registers(32)    <= not(registers(31));                                                                              
                registers(33)    <= not(registers(32));                                                                              
                registers(34)    <= not(registers(33));                                                                              
                registers(35)    <= not(registers(34));                                                                              
                registers(36)    <= not(registers(35));                                                                              
                registers(37)    <= not(registers(36));                                                                              
                registers(38)    <= not(registers(37));                                                                              
                registers(39)    <= not(registers(38));                                                                              
                registers(40)    <= not(registers(39));                                                                              
                registers(41)    <= not(registers(40));                                                                              
                registers(42)    <= not(registers(41));                                                                              
                registers(43)    <= not(registers(42));                                                                              
                registers(44)    <= not(registers(43));                                                                              
                registers(45)    <= not(registers(44));                                                                              
                registers(46)    <= not(registers(45));                                                                              
                registers(47)    <= not(registers(46));                                                                              
                registers(48)    <= not(registers(47));                                                                              
                registers(49)    <= not(registers(48));                                                                              
                registers(50)    <= not(registers(49));                                                                              
                registers(51)    <= not(registers(50));                                                                              
                registers(52)    <= not(registers(51));                                                                              
                registers(53)    <= not(registers(52));                                                                              
                registers(54)    <= not(registers(53));                                                                              
                registers(55)    <= not(registers(54));                                                                              
                registers(56)    <= not(registers(55));                                                                              
                registers(57)    <= not(registers(56));                                                                              
                registers(58)    <= not(registers(57));                                                                              
                registers(59)    <= not(registers(58));                                                                              
                registers(60)    <= not(registers(59));                                                                              
                registers(61)    <= not(registers(60));                                                                              
                registers(62)    <= not(registers(61));                                                                              
                registers(63)    <= not(registers(62));                                                                              
                registers(64)    <= not(registers(63));                                                                              
                registers(65)    <= not(registers(64));                                                                              
                registers(66)    <= not(registers(65));                                                                              
                registers(67)    <= not(registers(66));                                                                              
                registers(68)    <= not(registers(67));                                                                              
                registers(69)    <= not(registers(68));                                                                              
                registers(70)    <= not(registers(69));                                                                              
                registers(71)    <= not(registers(70));                                                                              
                registers(72)    <= not(registers(71));                                                                              
                registers(73)    <= not(registers(72));                                                                              
                registers(74)    <= not(registers(73));                                                                              
                registers(75)    <= not(registers(74));                                                                              
                registers(76)    <= not(registers(75));                                                                              
                registers(77)    <= not(registers(76));                                                                              
                registers(78)    <= not(registers(77));                                                                              
                registers(79)    <= not(registers(78));                                                                              
                registers(80)    <= not(registers(79));                                                                              
                registers(81)    <= not(registers(80));                                                                              
                registers(82)    <= not(registers(81));                                                                              
                registers(83)    <= not(registers(82));                                                                              
                registers(84)    <= not(registers(83));                                                                              
                registers(85)    <= not(registers(84));                                                                              
                registers(86)    <= not(registers(85));                                                                              
                registers(87)    <= not(registers(86));                                                                              
                registers(88)    <= not(registers(87));                                                                              
                registers(89)    <= not(registers(88));                                                                              
                registers(90)    <= not(registers(89));                                                                              
                registers(91)    <= not(registers(90));                                                                              
                registers(92)    <= not(registers(91));                                                                              
                registers(93)    <= not(registers(92));                                                                              
                registers(94)    <= not(registers(93));                                                                              
                registers(95)    <= not(registers(94));                                                                              
                registers(96)    <= not(registers(95));                                                                              
                registers(97)    <= not(registers(96));                                                                              
                registers(98)    <= not(registers(97));                                                                              
                registers(99)    <= not(registers(98));                                                                              
                registers(100)    <= not(registers(99));                                                                              
                registers(101)    <= not(registers(100));                                                                              
                registers(102)    <= not(registers(101));                                                                              
                registers(103)    <= not(registers(102));                                                                              
                registers(104)    <= not(registers(103));                                                                              
                registers(105)    <= not(registers(104));                                                                              
                registers(106)    <= not(registers(105));                                                                              
                registers(107)    <= not(registers(106));                                                                              
                registers(108)    <= not(registers(107));                                                                              
                registers(109)    <= not(registers(108));                                                                              
                registers(110)    <= not(registers(109));                                                                              
                registers(111)    <= not(registers(110));                                                                              
                registers(112)    <= not(registers(111));                                                                              
                registers(113)    <= not(registers(112));                                                                              
                registers(114)    <= not(registers(113));                                                                              
                registers(115)    <= not(registers(114));                                                                              
                registers(116)    <= not(registers(115));                                                                              
                registers(117)    <= not(registers(116));                                                                              
                registers(118)    <= not(registers(117));                                                                              
                registers(119)    <= not(registers(118));                                                                              
                registers(120)    <= not(registers(119));                                                                              
                registers(121)    <= not(registers(120));                                                                              
                registers(122)    <= not(registers(121));                                                                              
                registers(123)    <= not(registers(122));                                                                              
                registers(124)    <= not(registers(123));                                                                              
                registers(125)    <= not(registers(124));                                                                              
                registers(126)    <= not(registers(125));                                                                              
                registers(127)    <= not(registers(126));                                                                              
                registers(128)    <= not(registers(127));                                                                              
                registers(129)    <= not(registers(128));                                                                              
                registers(130)    <= not(registers(129));                                                                              
                registers(131)    <= not(registers(130));                                                                              
                registers(132)    <= not(registers(131));                                                                              
                registers(133)    <= not(registers(132));                                                                              
                registers(134)    <= not(registers(133));                                                                              
                registers(135)    <= not(registers(134));                                                                              
                registers(136)    <= not(registers(135));                                                                              
                registers(137)    <= not(registers(136));                                                                              
                registers(138)    <= not(registers(137));                                                                              
                registers(139)    <= not(registers(138));                                                                              
                registers(140)    <= not(registers(139));                                                                              
                registers(141)    <= not(registers(140));                                                                              
                registers(142)    <= not(registers(141));                                                                              
                registers(143)    <= not(registers(142));                                                                              
                registers(144)    <= not(registers(143));                                                                              
                registers(145)    <= not(registers(144));                                                                              
                registers(146)    <= not(registers(145));                                                                              
                registers(147)    <= not(registers(146));                                                                              
                registers(148)    <= not(registers(147));                                                                              
                registers(149)    <= not(registers(148));                                                                              
                registers(150)    <= not(registers(149));                                                                              
                registers(151)    <= not(registers(150));                                                                              
                registers(152)    <= not(registers(151));                                                                              
                registers(153)    <= not(registers(152));                                                                              
                registers(154)    <= not(registers(153));                                                                              
                registers(155)    <= not(registers(154));                                                                              
                registers(156)    <= not(registers(155));                                                                              
                registers(157)    <= not(registers(156));                                                                              
                registers(158)    <= not(registers(157));                                                                              
                registers(159)    <= not(registers(158));                                                                              
                registers(160)    <= not(registers(159));                                                                              
                registers(161)    <= not(registers(160));                                                                              
                registers(162)    <= not(registers(161));                                                                              
                registers(163)    <= not(registers(162));                                                                              
                registers(164)    <= not(registers(163));                                                                              
                registers(165)    <= not(registers(164));                                                                              
                registers(166)    <= not(registers(165));                                                                              
                registers(167)    <= not(registers(166));                                                                              
                registers(168)    <= not(registers(167));                                                                              
                registers(169)    <= not(registers(168));                                                                              
                registers(170)    <= not(registers(169));                                                                              
                registers(171)    <= not(registers(170));                                                                              
                registers(172)    <= not(registers(171));                                                                              
                registers(173)    <= not(registers(172));                                                                              
                registers(174)    <= not(registers(173));                                                                              
                registers(175)    <= not(registers(174));                                                                              
                registers(176)    <= not(registers(175));                                                                              
                registers(177)    <= not(registers(176));                                                                              
                registers(178)    <= not(registers(177));                                                                              
                registers(179)    <= not(registers(178));                                                                              
                registers(180)    <= not(registers(179));                                                                              
                registers(181)    <= not(registers(180));                                                                              
                registers(182)    <= not(registers(181));                                                                              
                registers(183)    <= not(registers(182));                                                                              
                registers(184)    <= not(registers(183));                                                                              
                registers(185)    <= not(registers(184));                                                                              
                registers(186)    <= not(registers(185));                                                                              
                registers(187)    <= not(registers(186));                                                                              
                registers(188)    <= not(registers(187));                                                                              
                registers(189)    <= not(registers(188));                                                                              
                registers(190)    <= not(registers(189));                                                                              
                registers(191)    <= not(registers(190));                                                                              
                registers(192)    <= not(registers(191));                                                                              
                registers(193)    <= not(registers(192));                                                                              
                registers(194)    <= not(registers(193));                                                                              
                registers(195)    <= not(registers(194));                                                                              
                registers(196)    <= not(registers(195));                                                                              
                registers(197)    <= not(registers(196));                                                                              
                registers(198)    <= not(registers(197));                                                                              
                registers(199)    <= not(registers(198));                                                                              
                registers(200)    <= not(registers(199));                                                                              
                registers(201)    <= not(registers(200));                                                                              
                registers(202)    <= not(registers(201));                                                                              
                registers(203)    <= not(registers(202));                                                                              
                registers(204)    <= not(registers(203));                                                                              
                registers(205)    <= not(registers(204));                                                                              
                registers(206)    <= not(registers(205));                                                                              
                registers(207)    <= not(registers(206));                                                                              
                registers(208)    <= not(registers(207));                                                                              
                registers(209)    <= not(registers(208));                                                                              
                registers(210)    <= not(registers(209));                                                                              
                registers(211)    <= not(registers(210));                                                                              
                registers(212)    <= not(registers(211));                                                                              
                registers(213)    <= not(registers(212));                                                                              
                registers(214)    <= not(registers(213));                                                                              
                registers(215)    <= not(registers(214));                                                                              
                registers(216)    <= not(registers(215));                                                                              
                registers(217)    <= not(registers(216));                                                                              
                registers(218)    <= not(registers(217));                                                                              
                registers(219)    <= not(registers(218));                                                                              
                registers(220)    <= not(registers(219));                                                                              
                registers(221)    <= not(registers(220));                                                                              
                registers(222)    <= not(registers(221));                                                                              
                registers(223)    <= not(registers(222));                                                                              
                registers(224)    <= not(registers(223));                                                                              
                registers(225)    <= not(registers(224));                                                                              
                registers(226)    <= not(registers(225));                                                                              
                registers(227)    <= not(registers(226));                                                                              
                registers(228)    <= not(registers(227));                                                                              
                registers(229)    <= not(registers(228));                                                                              
                registers(230)    <= not(registers(229));                                                                              
                registers(231)    <= not(registers(230));                                                                              
                registers(232)    <= not(registers(231));                                                                              
                registers(233)    <= not(registers(232));                                                                              
                registers(234)    <= not(registers(233));                                                                              
                registers(235)    <= not(registers(234));                                                                              
                registers(236)    <= not(registers(235));                                                                              
                registers(237)    <= not(registers(236));                                                                              
                registers(238)    <= not(registers(237));                                                                              
                registers(239)    <= not(registers(238));                                                                              
                registers(240)    <= not(registers(239));                                                                              
                registers(241)    <= not(registers(240));                                                                              
                registers(242)    <= not(registers(241));                                                                              
                registers(243)    <= not(registers(242));                                                                              
                registers(244)    <= not(registers(243));                                                                              
                registers(245)    <= not(registers(244));                                                                              
                registers(246)    <= not(registers(245));                                                                              
                registers(247)    <= not(registers(246));                                                                              
                registers(248)    <= not(registers(247));                                                                              
                registers(249)    <= not(registers(248));                                                                              
                registers(250)    <= not(registers(249));                                                                              
                registers(251)    <= not(registers(250));                                                                              
                registers(252)    <= not(registers(251));                                                                              
                registers(253)    <= not(registers(252));                                                                              
                registers(254)    <= not(registers(253));                                                                              
                registers(255)    <= not(registers(254));                                                                              
                registers(256)    <= not(registers(255));                                                                              
                registers(257)    <= not(registers(256));                                                                              
                registers(258)    <= not(registers(257));                                                                              
                registers(259)    <= not(registers(258));                                                                              
                registers(260)    <= not(registers(259));                                                                              
                registers(261)    <= not(registers(260));                                                                              
                registers(262)    <= not(registers(261));                                                                              
                registers(263)    <= not(registers(262));                                                                              
                registers(264)    <= not(registers(263));                                                                              
                registers(265)    <= not(registers(264));                                                                              
                registers(266)    <= not(registers(265));                                                                              
                registers(267)    <= not(registers(266));                                                                              
                registers(268)    <= not(registers(267));                                                                              
                registers(269)    <= not(registers(268));                                                                              
                registers(270)    <= not(registers(269));                                                                              
                registers(271)    <= not(registers(270));                                                                              
                registers(272)    <= not(registers(271));                                                                              
                registers(273)    <= not(registers(272));                                                                              
                registers(274)    <= not(registers(273));                                                                              
                registers(275)    <= not(registers(274));                                                                              
                registers(276)    <= not(registers(275));                                                                              
                registers(277)    <= not(registers(276));                                                                              
                registers(278)    <= not(registers(277));                                                                              
                registers(279)    <= not(registers(278));                                                                              
                registers(280)    <= not(registers(279));                                                                              
                registers(281)    <= not(registers(280));                                                                              
                registers(282)    <= not(registers(281));                                                                              
                registers(283)    <= not(registers(282));                                                                              
                registers(284)    <= not(registers(283));                                                                              
                registers(285)    <= not(registers(284));                                                                              
                registers(286)    <= not(registers(285));                                                                              
                registers(287)    <= not(registers(286));                                                                              
                registers(288)    <= not(registers(287));                                                                              
                registers(289)    <= not(registers(288));                                                                              
                registers(290)    <= not(registers(289));                                                                              
                registers(291)    <= not(registers(290));                                                                              
                registers(292)    <= not(registers(291));                                                                              
                registers(293)    <= not(registers(292));                                                                              
                registers(294)    <= not(registers(293));                                                                              
                registers(295)    <= not(registers(294));                                                                              
                registers(296)    <= not(registers(295));                                                                              
                registers(297)    <= not(registers(296));                                                                              
                registers(298)    <= not(registers(297));                                                                              
                registers(299)    <= not(registers(298));                                                                              
                registers(300)    <= not(registers(299));                                                                              
                registers(301)    <= not(registers(300));                                                                              
                registers(302)    <= not(registers(301));                                                                              
                registers(303)    <= not(registers(302));                                                                              
                registers(304)    <= not(registers(303));                                                                              
                registers(305)    <= not(registers(304));                                                                              
                registers(306)    <= not(registers(305));                                                                              
                registers(307)    <= not(registers(306));                                                                              
                registers(308)    <= not(registers(307));                                                                              
                registers(309)    <= not(registers(308));                                                                              
                registers(310)    <= not(registers(309));                                                                              
                registers(311)    <= not(registers(310));                                                                              
                registers(312)    <= not(registers(311));                                                                              
                registers(313)    <= not(registers(312));                                                                              
                registers(314)    <= not(registers(313));                                                                              
                registers(315)    <= not(registers(314));                                                                              
                registers(316)    <= not(registers(315));                                                                              
                registers(317)    <= not(registers(316));                                                                              
                registers(318)    <= not(registers(317));                                                                              
                registers(319)    <= not(registers(318));                                                                              
                registers(320)    <= not(registers(319));                                                                              
                registers(321)    <= not(registers(320));                                                                              
                registers(322)    <= not(registers(321));                                                                              
                registers(323)    <= not(registers(322));                                                                              
                registers(324)    <= not(registers(323));                                                                              
                registers(325)    <= not(registers(324));                                                                              
                registers(326)    <= not(registers(325));                                                                              
                registers(327)    <= not(registers(326));                                                                              
                registers(328)    <= not(registers(327));                                                                              
                registers(329)    <= not(registers(328));                                                                              
                registers(330)    <= not(registers(329));                                                                              
                registers(331)    <= not(registers(330));                                                                              
                registers(332)    <= not(registers(331));                                                                              
                registers(333)    <= not(registers(332));                                                                              
                registers(334)    <= not(registers(333));                                                                              
                registers(335)    <= not(registers(334));                                                                              
                registers(336)    <= not(registers(335));                                                                              
                registers(337)    <= not(registers(336));                                                                              
                registers(338)    <= not(registers(337));                                                                              
                registers(339)    <= not(registers(338));                                                                              
                registers(340)    <= not(registers(339));                                                                              
                registers(341)    <= not(registers(340));                                                                              
                registers(342)    <= not(registers(341));                                                                              
                registers(343)    <= not(registers(342));                                                                              
                registers(344)    <= not(registers(343));                                                                              
                registers(345)    <= not(registers(344));                                                                              
                registers(346)    <= not(registers(345));                                                                              
                registers(347)    <= not(registers(346));                                                                              
                registers(348)    <= not(registers(347));                                                                              
                registers(349)    <= not(registers(348));                                                                              
                registers(350)    <= not(registers(349));                                                                              
                registers(351)    <= not(registers(350));                                                                              
                registers(352)    <= not(registers(351));                                                                              
                registers(353)    <= not(registers(352));                                                                              
                registers(354)    <= not(registers(353));                                                                              
                registers(355)    <= not(registers(354));                                                                              
                registers(356)    <= not(registers(355));                                                                              
                registers(357)    <= not(registers(356));                                                                              
                registers(358)    <= not(registers(357));                                                                              
                registers(359)    <= not(registers(358));                                                                              
                registers(360)    <= not(registers(359));                                                                              
                registers(361)    <= not(registers(360));                                                                              
                registers(362)    <= not(registers(361));                                                                              
                registers(363)    <= not(registers(362));                                                                              
                registers(364)    <= not(registers(363));                                                                              
                registers(365)    <= not(registers(364));                                                                              
                registers(366)    <= not(registers(365));                                                                              
                registers(367)    <= not(registers(366));                                                                              
                registers(368)    <= not(registers(367));                                                                              
                registers(369)    <= not(registers(368));                                                                              
                registers(370)    <= not(registers(369));                                                                              
                registers(371)    <= not(registers(370));                                                                              
                registers(372)    <= not(registers(371));                                                                              
                registers(373)    <= not(registers(372));                                                                              
                registers(374)    <= not(registers(373));                                                                              
                registers(375)    <= not(registers(374));                                                                              
                registers(376)    <= not(registers(375));                                                                              
                registers(377)    <= not(registers(376));                                                                              
                registers(378)    <= not(registers(377));                                                                              
                registers(379)    <= not(registers(378));                                                                              
                registers(380)    <= not(registers(379));                                                                              
                registers(381)    <= not(registers(380));                                                                              
                registers(382)    <= not(registers(381));                                                                              
                registers(383)    <= not(registers(382));                                                                              
                registers(384)    <= not(registers(383));                                                                              
                registers(385)    <= not(registers(384));                                                                              
                registers(386)    <= not(registers(385));                                                                              
                registers(387)    <= not(registers(386));                                                                              
                registers(388)    <= not(registers(387));                                                                              
                registers(389)    <= not(registers(388));                                                                              
                registers(390)    <= not(registers(389));                                                                              
                registers(391)    <= not(registers(390));                                                                              
                registers(392)    <= not(registers(391));                                                                              
                registers(393)    <= not(registers(392));                                                                              
                registers(394)    <= not(registers(393));                                                                              
                registers(395)    <= not(registers(394));                                                                              
                registers(396)    <= not(registers(395));                                                                              
                registers(397)    <= not(registers(396));                                                                              
                registers(398)    <= not(registers(397));                                                                              
                registers(399)    <= not(registers(398));                                                                              
                registers(400)    <= not(registers(399));                                                                              
                registers(401)    <= not(registers(400));                                                                              
                registers(402)    <= not(registers(401));                                                                              
                registers(403)    <= not(registers(402));                                                                              
                registers(404)    <= not(registers(403));                                                                              
                registers(405)    <= not(registers(404));                                                                              
                registers(406)    <= not(registers(405));                                                                              
                registers(407)    <= not(registers(406));                                                                              
                registers(408)    <= not(registers(407));                                                                              
                registers(409)    <= not(registers(408));                                                                              
                registers(410)    <= not(registers(409));                                                                              
                registers(411)    <= not(registers(410));                                                                              
                registers(412)    <= not(registers(411));                                                                              
                registers(413)    <= not(registers(412));                                                                              
                registers(414)    <= not(registers(413));                                                                              
                registers(415)    <= not(registers(414));                                                                              
                registers(416)    <= not(registers(415));                                                                              
                registers(417)    <= not(registers(416));                                                                              
                registers(418)    <= not(registers(417));                                                                              
                registers(419)    <= not(registers(418));                                                                              
                registers(420)    <= not(registers(419));                                                                              
                registers(421)    <= not(registers(420));                                                                              
                registers(422)    <= not(registers(421));                                                                              
                registers(423)    <= not(registers(422));                                                                              
                registers(424)    <= not(registers(423));                                                                              
                registers(425)    <= not(registers(424));                                                                              
                registers(426)    <= not(registers(425));                                                                              
                registers(427)    <= not(registers(426));                                                                              
                registers(428)    <= not(registers(427));                                                                              
                registers(429)    <= not(registers(428));                                                                              
                registers(430)    <= not(registers(429));                                                                              
                registers(431)    <= not(registers(430));                                                                              
                registers(432)    <= not(registers(431));                                                                              
                registers(433)    <= not(registers(432));                                                                              
                registers(434)    <= not(registers(433));                                                                              
                registers(435)    <= not(registers(434));                                                                              
                registers(436)    <= not(registers(435));                                                                              
                registers(437)    <= not(registers(436));                                                                              
                registers(438)    <= not(registers(437));                                                                              
                registers(439)    <= not(registers(438));                                                                              
                registers(440)    <= not(registers(439));                                                                              
                registers(441)    <= not(registers(440));                                                                              
                registers(442)    <= not(registers(441));                                                                              
                registers(443)    <= not(registers(442));                                                                              
                registers(444)    <= not(registers(443));                                                                              
                registers(445)    <= not(registers(444));                                                                              
                registers(446)    <= not(registers(445));                                                                              
                registers(447)    <= not(registers(446));                                                                              
                registers(448)    <= not(registers(447));                                                                              
                registers(449)    <= not(registers(448));                                                                              
                registers(450)    <= not(registers(449));                                                                              
                registers(451)    <= not(registers(450));                                                                              
                registers(452)    <= not(registers(451));                                                                              
                registers(453)    <= not(registers(452));                                                                              
                registers(454)    <= not(registers(453));                                                                              
                registers(455)    <= not(registers(454));                                                                              
                registers(456)    <= not(registers(455));                                                                              
                registers(457)    <= not(registers(456));                                                                              
                registers(458)    <= not(registers(457));                                                                              
                registers(459)    <= not(registers(458));                                                                              
                registers(460)    <= not(registers(459));                                                                              
                registers(461)    <= not(registers(460));                                                                              
                registers(462)    <= not(registers(461));                                                                              
                registers(463)    <= not(registers(462));                                                                              
                registers(464)    <= not(registers(463));                                                                              
                registers(465)    <= not(registers(464));                                                                              
                registers(466)    <= not(registers(465));                                                                              
                registers(467)    <= not(registers(466));                                                                              
                registers(468)    <= not(registers(467));                                                                              
                registers(469)    <= not(registers(468));                                                                              
                registers(470)    <= not(registers(469));                                                                              
                registers(471)    <= not(registers(470));                                                                              
                registers(472)    <= not(registers(471));                                                                              
                registers(473)    <= not(registers(472));                                                                              
                registers(474)    <= not(registers(473));                                                                              
                registers(475)    <= not(registers(474));                                                                              
                registers(476)    <= not(registers(475));                                                                              
                registers(477)    <= not(registers(476));                                                                              
                registers(478)    <= not(registers(477));                                                                              
                registers(479)    <= not(registers(478));                                                                              
                registers(480)    <= not(registers(479));                                                                              
                registers(481)    <= not(registers(480));                                                                              
                registers(482)    <= not(registers(481));                                                                              
                registers(483)    <= not(registers(482));                                                                              
                registers(484)    <= not(registers(483));                                                                              
                registers(485)    <= not(registers(484));                                                                              
                registers(486)    <= not(registers(485));                                                                              
                registers(487)    <= not(registers(486));                                                                              
                registers(488)    <= not(registers(487));                                                                              
                registers(489)    <= not(registers(488));                                                                              
                registers(490)    <= not(registers(489));                                                                              
                registers(491)    <= not(registers(490));                                                                              
                registers(492)    <= not(registers(491));                                                                              
                registers(493)    <= not(registers(492));                                                                              
                registers(494)    <= not(registers(493));                                                                              
                registers(495)    <= not(registers(494));                                                                              
                registers(496)    <= not(registers(495));                                                                              
                registers(497)    <= not(registers(496));                                                                              
                registers(498)    <= not(registers(497));                                                                              
                registers(499)    <= not(registers(498));                                                                              
                registers(500)    <= not(registers(499));                                                                              
                registers(501)    <= not(registers(500));                                                                              
                registers(502)    <= not(registers(501));                                                                              
                registers(503)    <= not(registers(502));                                                                              
                registers(504)    <= not(registers(503));                                                                              
                registers(505)    <= not(registers(504));                                                                              
                registers(506)    <= not(registers(505));                                                                              
                registers(507)    <= not(registers(506));                                                                              
                registers(508)    <= not(registers(507));                                                                              
                registers(509)    <= not(registers(508));                                                                              
                registers(510)    <= not(registers(509));                                                                              
                registers(511)    <= not(registers(510));                                                                              
                registers(512)    <= not(registers(511));                                                                              
                registers(513)    <= not(registers(512));                                                                              
                registers(514)    <= not(registers(513));                                                                              
                registers(515)    <= not(registers(514));                                                                              
                registers(516)    <= not(registers(515));                                                                              
                registers(517)    <= not(registers(516));                                                                              
                registers(518)    <= not(registers(517));                                                                              
                registers(519)    <= not(registers(518));                                                                              
                registers(520)    <= not(registers(519));                                                                              
                registers(521)    <= not(registers(520));                                                                              
                registers(522)    <= not(registers(521));                                                                              
                registers(523)    <= not(registers(522));                                                                              
                registers(524)    <= not(registers(523));                                                                              
                registers(525)    <= not(registers(524));                                                                              
                registers(526)    <= not(registers(525));                                                                              
                registers(527)    <= not(registers(526));                                                                              
                registers(528)    <= not(registers(527));                                                                              
                registers(529)    <= not(registers(528));                                                                              
                registers(530)    <= not(registers(529));                                                                              
                registers(531)    <= not(registers(530));                                                                              
                registers(532)    <= not(registers(531));                                                                              
                registers(533)    <= not(registers(532));                                                                              
                registers(534)    <= not(registers(533));                                                                              
                registers(535)    <= not(registers(534));                                                                              
                registers(536)    <= not(registers(535));                                                                              
                registers(537)    <= not(registers(536));                                                                              
                registers(538)    <= not(registers(537));                                                                              
                registers(539)    <= not(registers(538));                                                                              
                registers(540)    <= not(registers(539));                                                                              
                registers(541)    <= not(registers(540));                                                                              
                registers(542)    <= not(registers(541));                                                                              
                registers(543)    <= not(registers(542));                                                                              
                registers(544)    <= not(registers(543));                                                                              
                registers(545)    <= not(registers(544));                                                                              
                registers(546)    <= not(registers(545));                                                                              
                registers(547)    <= not(registers(546));                                                                              
                registers(548)    <= not(registers(547));                                                                              
                registers(549)    <= not(registers(548));                                                                              
                registers(550)    <= not(registers(549));                                                                              
                registers(551)    <= not(registers(550));                                                                              
                registers(552)    <= not(registers(551));                                                                              
                registers(553)    <= not(registers(552));                                                                              
                registers(554)    <= not(registers(553));                                                                              
                registers(555)    <= not(registers(554));                                                                              
                registers(556)    <= not(registers(555));                                                                              
                registers(557)    <= not(registers(556));                                                                              
                registers(558)    <= not(registers(557));                                                                              
                registers(559)    <= not(registers(558));                                                                              
                registers(560)    <= not(registers(559));                                                                              
                registers(561)    <= not(registers(560));                                                                              
                registers(562)    <= not(registers(561));                                                                              
                registers(563)    <= not(registers(562));                                                                              
                registers(564)    <= not(registers(563));                                                                              
                registers(565)    <= not(registers(564));                                                                              
                registers(566)    <= not(registers(565));                                                                              
                registers(567)    <= not(registers(566));                                                                              
                registers(568)    <= not(registers(567));                                                                              
                registers(569)    <= not(registers(568));                                                                              
                registers(570)    <= not(registers(569));                                                                              
                registers(571)    <= not(registers(570));                                                                              
                registers(572)    <= not(registers(571));                                                                              
                registers(573)    <= not(registers(572));                                                                              
                registers(574)    <= not(registers(573));                                                                              
                registers(575)    <= not(registers(574));                                                                              
                registers(576)    <= not(registers(575));                                                                              
                registers(577)    <= not(registers(576));                                                                              
                registers(578)    <= not(registers(577));                                                                              
                registers(579)    <= not(registers(578));                                                                              
                registers(580)    <= not(registers(579));                                                                              
                registers(581)    <= not(registers(580));                                                                              
                registers(582)    <= not(registers(581));                                                                              
                registers(583)    <= not(registers(582));                                                                              
                registers(584)    <= not(registers(583));                                                                              
                registers(585)    <= not(registers(584));                                                                              
                registers(586)    <= not(registers(585));                                                                              
                registers(587)    <= not(registers(586));                                                                              
                registers(588)    <= not(registers(587));                                                                              
                registers(589)    <= not(registers(588));                                                                              
                registers(590)    <= not(registers(589));                                                                              
                registers(591)    <= not(registers(590));                                                                              
                registers(592)    <= not(registers(591));                                                                              
                registers(593)    <= not(registers(592));                                                                              
                registers(594)    <= not(registers(593));                                                                              
                registers(595)    <= not(registers(594));                                                                              
                registers(596)    <= not(registers(595));                                                                              
                registers(597)    <= not(registers(596));                                                                              
                registers(598)    <= not(registers(597));                                                                              
                registers(599)    <= not(registers(598));                                                                              
                registers(600)    <= not(registers(599));                                                                              
                registers(601)    <= not(registers(600));                                                                              
                registers(602)    <= not(registers(601));                                                                              
                registers(603)    <= not(registers(602));                                                                              
                registers(604)    <= not(registers(603));                                                                              
                registers(605)    <= not(registers(604));                                                                              
                registers(606)    <= not(registers(605));                                                                              
                registers(607)    <= not(registers(606));                                                                              
                registers(608)    <= not(registers(607));                                                                              
                registers(609)    <= not(registers(608));                                                                              
                registers(610)    <= not(registers(609));                                                                              
                registers(611)    <= not(registers(610));                                                                              
                registers(612)    <= not(registers(611));                                                                              
                registers(613)    <= not(registers(612));                                                                              
                registers(614)    <= not(registers(613));                                                                              
                registers(615)    <= not(registers(614));                                                                              
                registers(616)    <= not(registers(615));                                                                              
                registers(617)    <= not(registers(616));                                                                              
                registers(618)    <= not(registers(617));                                                                              
                registers(619)    <= not(registers(618));                                                                              
                registers(620)    <= not(registers(619));                                                                              
                registers(621)    <= not(registers(620));                                                                              
                registers(622)    <= not(registers(621));                                                                              
                registers(623)    <= not(registers(622));                                                                              
                registers(624)    <= not(registers(623));                                                                              
                registers(625)    <= not(registers(624));                                                                              
                registers(626)    <= not(registers(625));                                                                              
                registers(627)    <= not(registers(626));                                                                              
                registers(628)    <= not(registers(627));                                                                              
                registers(629)    <= not(registers(628));                                                                              
                registers(630)    <= not(registers(629));                                                                              
                registers(631)    <= not(registers(630));                                                                              
                registers(632)    <= not(registers(631));                                                                              
                registers(633)    <= not(registers(632));                                                                              
                registers(634)    <= not(registers(633));                                                                              
                registers(635)    <= not(registers(634));                                                                              
                registers(636)    <= not(registers(635));                                                                              
                registers(637)    <= not(registers(636));                                                                              
                registers(638)    <= not(registers(637));                                                                              
                registers(639)    <= not(registers(638));                                                                              
                registers(640)    <= not(registers(639));                                                                              
                registers(641)    <= not(registers(640));                                                                              
                registers(642)    <= not(registers(641));                                                                              
                registers(643)    <= not(registers(642));                                                                              
                registers(644)    <= not(registers(643));                                                                              
                registers(645)    <= not(registers(644));                                                                              
                registers(646)    <= not(registers(645));                                                                              
                registers(647)    <= not(registers(646));                                                                              
                registers(648)    <= not(registers(647));                                                                              
                registers(649)    <= not(registers(648));                                                                              
                registers(650)    <= not(registers(649));                                                                              
                registers(651)    <= not(registers(650));                                                                              
                registers(652)    <= not(registers(651));                                                                              
                registers(653)    <= not(registers(652));                                                                              
                registers(654)    <= not(registers(653));                                                                              
                registers(655)    <= not(registers(654));                                                                              
                registers(656)    <= not(registers(655));                                                                              
                registers(657)    <= not(registers(656));                                                                              
                registers(658)    <= not(registers(657));                                                                              
                registers(659)    <= not(registers(658));                                                                              
                registers(660)    <= not(registers(659));                                                                              
                registers(661)    <= not(registers(660));                                                                              
                registers(662)    <= not(registers(661));                                                                              
                registers(663)    <= not(registers(662));                                                                              
                registers(664)    <= not(registers(663));                                                                              
                registers(665)    <= not(registers(664));                                                                              
                registers(666)    <= not(registers(665));                                                                              
                registers(667)    <= not(registers(666));                                                                              
                registers(668)    <= not(registers(667));                                                                              
                registers(669)    <= not(registers(668));                                                                              
                registers(670)    <= not(registers(669));                                                                              
                registers(671)    <= not(registers(670));                                                                              
                registers(672)    <= not(registers(671));                                                                              
                registers(673)    <= not(registers(672));                                                                              
                registers(674)    <= not(registers(673));                                                                              
                registers(675)    <= not(registers(674));                                                                              
                registers(676)    <= not(registers(675));                                                                              
                registers(677)    <= not(registers(676));                                                                              
                registers(678)    <= not(registers(677));                                                                              
                registers(679)    <= not(registers(678));                                                                              
                registers(680)    <= not(registers(679));                                                                              
                registers(681)    <= not(registers(680));                                                                              
                registers(682)    <= not(registers(681));                                                                              
                registers(683)    <= not(registers(682));                                                                              
                registers(684)    <= not(registers(683));                                                                              
                registers(685)    <= not(registers(684));                                                                              
                registers(686)    <= not(registers(685));                                                                              
                registers(687)    <= not(registers(686));                                                                              
                registers(688)    <= not(registers(687));                                                                              
                registers(689)    <= not(registers(688));                                                                              
                registers(690)    <= not(registers(689));                                                                              
                registers(691)    <= not(registers(690));                                                                              
                registers(692)    <= not(registers(691));                                                                              
                registers(693)    <= not(registers(692));                                                                              
                registers(694)    <= not(registers(693));                                                                              
                registers(695)    <= not(registers(694));                                                                              
                registers(696)    <= not(registers(695));                                                                              
                registers(697)    <= not(registers(696));                                                                              
                registers(698)    <= not(registers(697));                                                                              
                registers(699)    <= not(registers(698));                                                                              
                registers(700)    <= not(registers(699));                                                                              
                registers(701)    <= not(registers(700));                                                                              
                registers(702)    <= not(registers(701));                                                                              
                registers(703)    <= not(registers(702));                                                                              
                registers(704)    <= not(registers(703));                                                                              
                registers(705)    <= not(registers(704));                                                                              
                registers(706)    <= not(registers(705));                                                                              
                registers(707)    <= not(registers(706));                                                                              
                registers(708)    <= not(registers(707));                                                                              
                registers(709)    <= not(registers(708));                                                                              
                registers(710)    <= not(registers(709));                                                                              
                registers(711)    <= not(registers(710));                                                                              
                registers(712)    <= not(registers(711));                                                                              
                registers(713)    <= not(registers(712));                                                                              
                registers(714)    <= not(registers(713));                                                                              
                registers(715)    <= not(registers(714));                                                                              
                registers(716)    <= not(registers(715));                                                                              
                registers(717)    <= not(registers(716));                                                                              
                registers(718)    <= not(registers(717));                                                                              
                registers(719)    <= not(registers(718));                                                                              
                registers(720)    <= not(registers(719));                                                                              
                registers(721)    <= not(registers(720));                                                                              
                registers(722)    <= not(registers(721));                                                                              
                registers(723)    <= not(registers(722));                                                                              
                registers(724)    <= not(registers(723));                                                                              
                registers(725)    <= not(registers(724));                                                                              
                registers(726)    <= not(registers(725));                                                                              
                registers(727)    <= not(registers(726));                                                                              
                registers(728)    <= not(registers(727));                                                                              
                registers(729)    <= not(registers(728));                                                                              
                registers(730)    <= not(registers(729));                                                                              
                registers(731)    <= not(registers(730));                                                                              
                registers(732)    <= not(registers(731));                                                                              
                registers(733)    <= not(registers(732));                                                                              
                registers(734)    <= not(registers(733));                                                                              
                registers(735)    <= not(registers(734));                                                                              
                registers(736)    <= not(registers(735));                                                                              
                registers(737)    <= not(registers(736));                                                                              
                registers(738)    <= not(registers(737));                                                                              
                registers(739)    <= not(registers(738));                                                                              
                registers(740)    <= not(registers(739));                                                                              
                registers(741)    <= not(registers(740));                                                                              
                registers(742)    <= not(registers(741));                                                                              
                registers(743)    <= not(registers(742));                                                                              
                registers(744)    <= not(registers(743));                                                                              
                registers(745)    <= not(registers(744));                                                                              
                registers(746)    <= not(registers(745));                                                                              
                registers(747)    <= not(registers(746));                                                                              
                registers(748)    <= not(registers(747));                                                                              
                registers(749)    <= not(registers(748));                                                                              
                registers(750)    <= not(registers(749));                                                                              
                registers(751)    <= not(registers(750));                                                                              
                registers(752)    <= not(registers(751));                                                                              
                registers(753)    <= not(registers(752));                                                                              
                registers(754)    <= not(registers(753));                                                                              
                registers(755)    <= not(registers(754));                                                                              
                registers(756)    <= not(registers(755));                                                                              
                registers(757)    <= not(registers(756));                                                                              
                registers(758)    <= not(registers(757));                                                                              
                registers(759)    <= not(registers(758));                                                                              
                registers(760)    <= not(registers(759));                                                                              
                registers(761)    <= not(registers(760));                                                                              
                registers(762)    <= not(registers(761));                                                                              
                registers(763)    <= not(registers(762));                                                                              
                registers(764)    <= not(registers(763));                                                                              
                registers(765)    <= not(registers(764));                                                                              
                registers(766)    <= not(registers(765));                                                                              
                registers(767)    <= not(registers(766));                                                                              
                registers(768)    <= not(registers(767));                                                                              
                registers(769)    <= not(registers(768));                                                                              
                registers(770)    <= not(registers(769));                                                                              
                registers(771)    <= not(registers(770));                                                                              
                registers(772)    <= not(registers(771));                                                                              
                registers(773)    <= not(registers(772));                                                                              
                registers(774)    <= not(registers(773));                                                                              
                registers(775)    <= not(registers(774));                                                                              
                registers(776)    <= not(registers(775));                                                                              
                registers(777)    <= not(registers(776));                                                                              
                registers(778)    <= not(registers(777));                                                                              
                registers(779)    <= not(registers(778));                                                                              
                registers(780)    <= not(registers(779));                                                                              
                registers(781)    <= not(registers(780));                                                                              
                registers(782)    <= not(registers(781));                                                                              
                registers(783)    <= not(registers(782));                                                                              
                registers(784)    <= not(registers(783));                                                                              
                registers(785)    <= not(registers(784));                                                                              
                registers(786)    <= not(registers(785));                                                                              
                registers(787)    <= not(registers(786));                                                                              
                registers(788)    <= not(registers(787));                                                                              
                registers(789)    <= not(registers(788));                                                                              
                registers(790)    <= not(registers(789));                                                                              
                registers(791)    <= not(registers(790));                                                                              
                registers(792)    <= not(registers(791));                                                                              
                registers(793)    <= not(registers(792));                                                                              
                registers(794)    <= not(registers(793));                                                                              
                registers(795)    <= not(registers(794));                                                                              
                registers(796)    <= not(registers(795));                                                                              
                registers(797)    <= not(registers(796));                                                                              
                registers(798)    <= not(registers(797));                                                                              
                registers(799)    <= not(registers(798));                                                                              
                registers(800)    <= not(registers(799));                                                                              
                registers(801)    <= not(registers(800));                                                                              
                registers(802)    <= not(registers(801));                                                                              
                registers(803)    <= not(registers(802));                                                                              
                registers(804)    <= not(registers(803));                                                                              
                registers(805)    <= not(registers(804));                                                                              
                registers(806)    <= not(registers(805));                                                                              
                registers(807)    <= not(registers(806));                                                                              
                registers(808)    <= not(registers(807));                                                                              
                registers(809)    <= not(registers(808));                                                                              
                registers(810)    <= not(registers(809));                                                                              
                registers(811)    <= not(registers(810));                                                                              
                registers(812)    <= not(registers(811));                                                                              
                registers(813)    <= not(registers(812));                                                                              
                registers(814)    <= not(registers(813));                                                                              
                registers(815)    <= not(registers(814));                                                                              
                registers(816)    <= not(registers(815));                                                                              
                registers(817)    <= not(registers(816));                                                                              
                registers(818)    <= not(registers(817));                                                                              
                registers(819)    <= not(registers(818));                                                                              
                registers(820)    <= not(registers(819));                                                                              
                registers(821)    <= not(registers(820));                                                                              
                registers(822)    <= not(registers(821));                                                                              
                registers(823)    <= not(registers(822));                                                                              
                registers(824)    <= not(registers(823));                                                                              
                registers(825)    <= not(registers(824));                                                                              
                registers(826)    <= not(registers(825));                                                                              
                registers(827)    <= not(registers(826));                                                                              
                registers(828)    <= not(registers(827));                                                                              
                registers(829)    <= not(registers(828));                                                                              
                registers(830)    <= not(registers(829));                                                                              
                registers(831)    <= not(registers(830));                                                                              
                registers(832)    <= not(registers(831));                                                                              
                registers(833)    <= not(registers(832));                                                                              
                registers(834)    <= not(registers(833));                                                                              
                registers(835)    <= not(registers(834));                                                                              
                registers(836)    <= not(registers(835));                                                                              
                registers(837)    <= not(registers(836));                                                                              
                registers(838)    <= not(registers(837));                                                                              
                registers(839)    <= not(registers(838));                                                                              
                registers(840)    <= not(registers(839));                                                                              
                registers(841)    <= not(registers(840));                                                                              
                registers(842)    <= not(registers(841));                                                                              
                registers(843)    <= not(registers(842));                                                                              
                registers(844)    <= not(registers(843));                                                                              
                registers(845)    <= not(registers(844));                                                                              
                registers(846)    <= not(registers(845));                                                                              
                registers(847)    <= not(registers(846));                                                                              
                registers(848)    <= not(registers(847));                                                                              
                registers(849)    <= not(registers(848));                                                                              
                registers(850)    <= not(registers(849));                                                                              
                registers(851)    <= not(registers(850));                                                                              
                registers(852)    <= not(registers(851));                                                                              
                registers(853)    <= not(registers(852));                                                                              
                registers(854)    <= not(registers(853));                                                                              
                registers(855)    <= not(registers(854));                                                                              
                registers(856)    <= not(registers(855));                                                                              
                registers(857)    <= not(registers(856));                                                                              
                registers(858)    <= not(registers(857));                                                                              
                registers(859)    <= not(registers(858));                                                                              
                registers(860)    <= not(registers(859));                                                                              
                registers(861)    <= not(registers(860));                                                                              
                registers(862)    <= not(registers(861));                                                                              
                registers(863)    <= not(registers(862));                                                                              
                registers(864)    <= not(registers(863));                                                                              
                registers(865)    <= not(registers(864));                                                                              
                registers(866)    <= not(registers(865));                                                                              
                registers(867)    <= not(registers(866));                                                                              
                registers(868)    <= not(registers(867));                                                                              
                registers(869)    <= not(registers(868));                                                                              
                registers(870)    <= not(registers(869));                                                                              
                registers(871)    <= not(registers(870));                                                                              
                registers(872)    <= not(registers(871));                                                                              
                registers(873)    <= not(registers(872));                                                                              
                registers(874)    <= not(registers(873));                                                                              
                registers(875)    <= not(registers(874));                                                                              
                registers(876)    <= not(registers(875));                                                                              
                registers(877)    <= not(registers(876));                                                                              
                registers(878)    <= not(registers(877));                                                                              
                registers(879)    <= not(registers(878));                                                                              
                registers(880)    <= not(registers(879));                                                                              
                registers(881)    <= not(registers(880));                                                                              
                registers(882)    <= not(registers(881));                                                                              
                registers(883)    <= not(registers(882));                                                                              
                registers(884)    <= not(registers(883));                                                                              
                registers(885)    <= not(registers(884));                                                                              
                registers(886)    <= not(registers(885));                                                                              
                registers(887)    <= not(registers(886));                                                                              
                registers(888)    <= not(registers(887));                                                                              
                registers(889)    <= not(registers(888));                                                                              
                registers(890)    <= not(registers(889));                                                                              
                registers(891)    <= not(registers(890));                                                                              
                registers(892)    <= not(registers(891));                                                                              
                registers(893)    <= not(registers(892));                                                                              
                registers(894)    <= not(registers(893));                                                                              
                registers(895)    <= not(registers(894));                                                                              
                registers(896)    <= not(registers(895));                                                                              
                registers(897)    <= not(registers(896));                                                                              
                registers(898)    <= not(registers(897));                                                                              
                registers(899)    <= not(registers(898));                                                                              
                registers(900)    <= not(registers(899));                                                                              
                registers(901)    <= not(registers(900));                                                                              
                registers(902)    <= not(registers(901));                                                                              
                registers(903)    <= not(registers(902));                                                                              
                registers(904)    <= not(registers(903));                                                                              
                registers(905)    <= not(registers(904));                                                                              
                registers(906)    <= not(registers(905));                                                                              
                registers(907)    <= not(registers(906));                                                                              
                registers(908)    <= not(registers(907));                                                                              
                registers(909)    <= not(registers(908));                                                                              
                registers(910)    <= not(registers(909));                                                                              
                registers(911)    <= not(registers(910));                                                                              
                registers(912)    <= not(registers(911));                                                                              
                registers(913)    <= not(registers(912));                                                                              
                registers(914)    <= not(registers(913));                                                                              
                registers(915)    <= not(registers(914));                                                                              
                registers(916)    <= not(registers(915));                                                                              
                registers(917)    <= not(registers(916));                                                                              
                registers(918)    <= not(registers(917));                                                                              
                registers(919)    <= not(registers(918));                                                                              
                registers(920)    <= not(registers(919));                                                                              
                registers(921)    <= not(registers(920));                                                                              
                registers(922)    <= not(registers(921));                                                                              
                registers(923)    <= not(registers(922));                                                                              
                registers(924)    <= not(registers(923));                                                                              
                registers(925)    <= not(registers(924));                                                                              
                registers(926)    <= not(registers(925));                                                                              
                registers(927)    <= not(registers(926));                                                                              
                registers(928)    <= not(registers(927));                                                                              
                registers(929)    <= not(registers(928));                                                                              
                registers(930)    <= not(registers(929));                                                                              
                registers(931)    <= not(registers(930));                                                                              
                registers(932)    <= not(registers(931));                                                                              
                registers(933)    <= not(registers(932));                                                                              
                registers(934)    <= not(registers(933));                                                                              
                registers(935)    <= not(registers(934));                                                                              
                registers(936)    <= not(registers(935));                                                                              
                registers(937)    <= not(registers(936));                                                                              
                registers(938)    <= not(registers(937));                                                                              
                registers(939)    <= not(registers(938));                                                                              
                registers(940)    <= not(registers(939));                                                                              
                registers(941)    <= not(registers(940));                                                                              
                registers(942)    <= not(registers(941));                                                                              
                registers(943)    <= not(registers(942));                                                                              
                registers(944)    <= not(registers(943));                                                                              
                registers(945)    <= not(registers(944));                                                                              
                registers(946)    <= not(registers(945));                                                                              
                registers(947)    <= not(registers(946));                                                                              
                registers(948)    <= not(registers(947));                                                                              
                registers(949)    <= not(registers(948));                                                                              
                registers(950)    <= not(registers(949));                                                                              
                registers(951)    <= not(registers(950));                                                                              
                registers(952)    <= not(registers(951));                                                                              
                registers(953)    <= not(registers(952));                                                                              
                registers(954)    <= not(registers(953));                                                                              
                registers(955)    <= not(registers(954));                                                                              
                registers(956)    <= not(registers(955));                                                                              
                registers(957)    <= not(registers(956));                                                                              
                registers(958)    <= not(registers(957));                                                                              
                registers(959)    <= not(registers(958));                                                                              
                registers(960)    <= not(registers(959));                                                                              
                registers(961)    <= not(registers(960));                                                                              
                registers(962)    <= not(registers(961));                                                                              
                registers(963)    <= not(registers(962));                                                                              
                registers(964)    <= not(registers(963));                                                                              
                registers(965)    <= not(registers(964));                                                                              
                registers(966)    <= not(registers(965));                                                                              
                registers(967)    <= not(registers(966));                                                                              
                registers(968)    <= not(registers(967));                                                                              
                registers(969)    <= not(registers(968));                                                                              
                registers(970)    <= not(registers(969));                                                                              
                registers(971)    <= not(registers(970));                                                                              
                registers(972)    <= not(registers(971));                                                                              
                registers(973)    <= not(registers(972));                                                                              
                registers(974)    <= not(registers(973));                                                                              
                registers(975)    <= not(registers(974));                                                                              
                registers(976)    <= not(registers(975));                                                                              
                registers(977)    <= not(registers(976));                                                                              
                registers(978)    <= not(registers(977));                                                                              
                registers(979)    <= not(registers(978));                                                                              
                registers(980)    <= not(registers(979));                                                                              
                registers(981)    <= not(registers(980));                                                                              
                registers(982)    <= not(registers(981));                                                                              
                registers(983)    <= not(registers(982));                                                                              
                registers(984)    <= not(registers(983));                                                                              
                registers(985)    <= not(registers(984));                                                                              
                registers(986)    <= not(registers(985));                                                                              
                registers(987)    <= not(registers(986));                                                                              
                registers(988)    <= not(registers(987));                                                                              
                registers(989)    <= not(registers(988));                                                                              
                registers(990)    <= not(registers(989));                                                                              
                registers(991)    <= not(registers(990));                                                                              
                registers(992)    <= not(registers(991));                                                                              
                registers(993)    <= not(registers(992));                                                                              
                registers(994)    <= not(registers(993));                                                                              
                registers(995)    <= not(registers(994));                                                                              
                registers(996)    <= not(registers(995));                                                                              
                registers(997)    <= not(registers(996));                                                                              
                registers(998)    <= not(registers(997));                                                                              
                registers(999)    <= not(registers(998));                                                                              
                                                                                                                                         
        end if;                                                                                                                          
    end process;                                                                                                                         
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Outputs                                                                                                                           
    ------------------------------------------                                                                                           
    process(clk)                                                                                                                         
    begin                                                                                                                                
                                                                                                                                         
        if rising_edge(clk) then                                                                                                         
                                                                                                                                         
            data_out(0) <= registers(nb_reg-4);                                                                                          
            data_out(1) <= registers(nb_reg-3);                                                                                          
            data_out(2) <= registers(nb_reg-2);                                                                                          
            data_out(3) <= registers(nb_reg-1);                                                                                          
                                                                                                                                         
        end if;                                                                                                                          
    end process;                                                                                                                         
                                                                                                                                         
end generate NO_MITIGATION;                                                                                                              
                                                                                                                                         
----------------------------------------------------------------------------------------------------------------------------             
--                                                                                                                                       
--                                                                                                                                       
--              Local TMR                                                                                                                
--                                                                                                                                       
--                                                                                                                                       
----------------------------------------------------------------------------------------------------------------------------             
                                                                                                                                         
LOCAL_TMR_MITIGATION: if USE_MITIGATION=1 generate                                                                                       
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Input                                                                                                                             
    ------------------------------------------                                                                                           
                                                                                                                                         
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Combinatiorial + Registers                                                                                                        
    ------------------------------------------                                                                                           
    process(clk)                                                                                                                         
    begin                                                                                                                                
                                                                                                                                         
        if rising_edge(clk) then                                                                                                         
                                                                                                                                         
                tmr_registers(0)(1)    <= not(local_tmr_voter(0));                                                                           
                tmr_registers(1)(1)    <= not(local_tmr_voter(0));                                                                           
                tmr_registers(2)(1)    <= not(local_tmr_voter(0));                                                                           
 
                tmr_registers(0)(2)    <= not(local_tmr_voter(1));                                                                           
                tmr_registers(1)(2)    <= not(local_tmr_voter(1));                                                                           
                tmr_registers(2)(2)    <= not(local_tmr_voter(1));                                                                           
 
                tmr_registers(0)(3)    <= not(local_tmr_voter(2));                                                                           
                tmr_registers(1)(3)    <= not(local_tmr_voter(2));                                                                           
                tmr_registers(2)(3)    <= not(local_tmr_voter(2));                                                                           
 
                tmr_registers(0)(4)    <= not(local_tmr_voter(3));                                                                           
                tmr_registers(1)(4)    <= not(local_tmr_voter(3));                                                                           
                tmr_registers(2)(4)    <= not(local_tmr_voter(3));                                                                           
 
                tmr_registers(0)(5)    <= not(local_tmr_voter(4));                                                                           
                tmr_registers(1)(5)    <= not(local_tmr_voter(4));                                                                           
                tmr_registers(2)(5)    <= not(local_tmr_voter(4));                                                                           
 
                tmr_registers(0)(6)    <= not(local_tmr_voter(5));                                                                           
                tmr_registers(1)(6)    <= not(local_tmr_voter(5));                                                                           
                tmr_registers(2)(6)    <= not(local_tmr_voter(5));                                                                           
 
                tmr_registers(0)(7)    <= not(local_tmr_voter(6));                                                                           
                tmr_registers(1)(7)    <= not(local_tmr_voter(6));                                                                           
                tmr_registers(2)(7)    <= not(local_tmr_voter(6));                                                                           
 
                tmr_registers(0)(8)    <= not(local_tmr_voter(7));                                                                           
                tmr_registers(1)(8)    <= not(local_tmr_voter(7));                                                                           
                tmr_registers(2)(8)    <= not(local_tmr_voter(7));                                                                           
 
                tmr_registers(0)(9)    <= not(local_tmr_voter(8));                                                                           
                tmr_registers(1)(9)    <= not(local_tmr_voter(8));                                                                           
                tmr_registers(2)(9)    <= not(local_tmr_voter(8));                                                                           
 
                tmr_registers(0)(10)    <= not(local_tmr_voter(9));                                                                           
                tmr_registers(1)(10)    <= not(local_tmr_voter(9));                                                                           
                tmr_registers(2)(10)    <= not(local_tmr_voter(9));                                                                           
 
                tmr_registers(0)(11)    <= not(local_tmr_voter(10));                                                                           
                tmr_registers(1)(11)    <= not(local_tmr_voter(10));                                                                           
                tmr_registers(2)(11)    <= not(local_tmr_voter(10));                                                                           
 
                tmr_registers(0)(12)    <= not(local_tmr_voter(11));                                                                           
                tmr_registers(1)(12)    <= not(local_tmr_voter(11));                                                                           
                tmr_registers(2)(12)    <= not(local_tmr_voter(11));                                                                           
 
                tmr_registers(0)(13)    <= not(local_tmr_voter(12));                                                                           
                tmr_registers(1)(13)    <= not(local_tmr_voter(12));                                                                           
                tmr_registers(2)(13)    <= not(local_tmr_voter(12));                                                                           
 
                tmr_registers(0)(14)    <= not(local_tmr_voter(13));                                                                           
                tmr_registers(1)(14)    <= not(local_tmr_voter(13));                                                                           
                tmr_registers(2)(14)    <= not(local_tmr_voter(13));                                                                           
 
                tmr_registers(0)(15)    <= not(local_tmr_voter(14));                                                                           
                tmr_registers(1)(15)    <= not(local_tmr_voter(14));                                                                           
                tmr_registers(2)(15)    <= not(local_tmr_voter(14));                                                                           
 
                tmr_registers(0)(16)    <= not(local_tmr_voter(15));                                                                           
                tmr_registers(1)(16)    <= not(local_tmr_voter(15));                                                                           
                tmr_registers(2)(16)    <= not(local_tmr_voter(15));                                                                           
 
                tmr_registers(0)(17)    <= not(local_tmr_voter(16));                                                                           
                tmr_registers(1)(17)    <= not(local_tmr_voter(16));                                                                           
                tmr_registers(2)(17)    <= not(local_tmr_voter(16));                                                                           
 
                tmr_registers(0)(18)    <= not(local_tmr_voter(17));                                                                           
                tmr_registers(1)(18)    <= not(local_tmr_voter(17));                                                                           
                tmr_registers(2)(18)    <= not(local_tmr_voter(17));                                                                           
 
                tmr_registers(0)(19)    <= not(local_tmr_voter(18));                                                                           
                tmr_registers(1)(19)    <= not(local_tmr_voter(18));                                                                           
                tmr_registers(2)(19)    <= not(local_tmr_voter(18));                                                                           
 
                tmr_registers(0)(20)    <= not(local_tmr_voter(19));                                                                           
                tmr_registers(1)(20)    <= not(local_tmr_voter(19));                                                                           
                tmr_registers(2)(20)    <= not(local_tmr_voter(19));                                                                           
 
                tmr_registers(0)(21)    <= not(local_tmr_voter(20));                                                                           
                tmr_registers(1)(21)    <= not(local_tmr_voter(20));                                                                           
                tmr_registers(2)(21)    <= not(local_tmr_voter(20));                                                                           
 
                tmr_registers(0)(22)    <= not(local_tmr_voter(21));                                                                           
                tmr_registers(1)(22)    <= not(local_tmr_voter(21));                                                                           
                tmr_registers(2)(22)    <= not(local_tmr_voter(21));                                                                           
 
                tmr_registers(0)(23)    <= not(local_tmr_voter(22));                                                                           
                tmr_registers(1)(23)    <= not(local_tmr_voter(22));                                                                           
                tmr_registers(2)(23)    <= not(local_tmr_voter(22));                                                                           
 
                tmr_registers(0)(24)    <= not(local_tmr_voter(23));                                                                           
                tmr_registers(1)(24)    <= not(local_tmr_voter(23));                                                                           
                tmr_registers(2)(24)    <= not(local_tmr_voter(23));                                                                           
 
                tmr_registers(0)(25)    <= not(local_tmr_voter(24));                                                                           
                tmr_registers(1)(25)    <= not(local_tmr_voter(24));                                                                           
                tmr_registers(2)(25)    <= not(local_tmr_voter(24));                                                                           
 
                tmr_registers(0)(26)    <= not(local_tmr_voter(25));                                                                           
                tmr_registers(1)(26)    <= not(local_tmr_voter(25));                                                                           
                tmr_registers(2)(26)    <= not(local_tmr_voter(25));                                                                           
 
                tmr_registers(0)(27)    <= not(local_tmr_voter(26));                                                                           
                tmr_registers(1)(27)    <= not(local_tmr_voter(26));                                                                           
                tmr_registers(2)(27)    <= not(local_tmr_voter(26));                                                                           
 
                tmr_registers(0)(28)    <= not(local_tmr_voter(27));                                                                           
                tmr_registers(1)(28)    <= not(local_tmr_voter(27));                                                                           
                tmr_registers(2)(28)    <= not(local_tmr_voter(27));                                                                           
 
                tmr_registers(0)(29)    <= not(local_tmr_voter(28));                                                                           
                tmr_registers(1)(29)    <= not(local_tmr_voter(28));                                                                           
                tmr_registers(2)(29)    <= not(local_tmr_voter(28));                                                                           
 
                tmr_registers(0)(30)    <= not(local_tmr_voter(29));                                                                           
                tmr_registers(1)(30)    <= not(local_tmr_voter(29));                                                                           
                tmr_registers(2)(30)    <= not(local_tmr_voter(29));                                                                           
 
                tmr_registers(0)(31)    <= not(local_tmr_voter(30));                                                                           
                tmr_registers(1)(31)    <= not(local_tmr_voter(30));                                                                           
                tmr_registers(2)(31)    <= not(local_tmr_voter(30));                                                                           
 
                tmr_registers(0)(32)    <= not(local_tmr_voter(31));                                                                           
                tmr_registers(1)(32)    <= not(local_tmr_voter(31));                                                                           
                tmr_registers(2)(32)    <= not(local_tmr_voter(31));                                                                           
 
                tmr_registers(0)(33)    <= not(local_tmr_voter(32));                                                                           
                tmr_registers(1)(33)    <= not(local_tmr_voter(32));                                                                           
                tmr_registers(2)(33)    <= not(local_tmr_voter(32));                                                                           
 
                tmr_registers(0)(34)    <= not(local_tmr_voter(33));                                                                           
                tmr_registers(1)(34)    <= not(local_tmr_voter(33));                                                                           
                tmr_registers(2)(34)    <= not(local_tmr_voter(33));                                                                           
 
                tmr_registers(0)(35)    <= not(local_tmr_voter(34));                                                                           
                tmr_registers(1)(35)    <= not(local_tmr_voter(34));                                                                           
                tmr_registers(2)(35)    <= not(local_tmr_voter(34));                                                                           
 
                tmr_registers(0)(36)    <= not(local_tmr_voter(35));                                                                           
                tmr_registers(1)(36)    <= not(local_tmr_voter(35));                                                                           
                tmr_registers(2)(36)    <= not(local_tmr_voter(35));                                                                           
 
                tmr_registers(0)(37)    <= not(local_tmr_voter(36));                                                                           
                tmr_registers(1)(37)    <= not(local_tmr_voter(36));                                                                           
                tmr_registers(2)(37)    <= not(local_tmr_voter(36));                                                                           
 
                tmr_registers(0)(38)    <= not(local_tmr_voter(37));                                                                           
                tmr_registers(1)(38)    <= not(local_tmr_voter(37));                                                                           
                tmr_registers(2)(38)    <= not(local_tmr_voter(37));                                                                           
 
                tmr_registers(0)(39)    <= not(local_tmr_voter(38));                                                                           
                tmr_registers(1)(39)    <= not(local_tmr_voter(38));                                                                           
                tmr_registers(2)(39)    <= not(local_tmr_voter(38));                                                                           
 
                tmr_registers(0)(40)    <= not(local_tmr_voter(39));                                                                           
                tmr_registers(1)(40)    <= not(local_tmr_voter(39));                                                                           
                tmr_registers(2)(40)    <= not(local_tmr_voter(39));                                                                           
 
                tmr_registers(0)(41)    <= not(local_tmr_voter(40));                                                                           
                tmr_registers(1)(41)    <= not(local_tmr_voter(40));                                                                           
                tmr_registers(2)(41)    <= not(local_tmr_voter(40));                                                                           
 
                tmr_registers(0)(42)    <= not(local_tmr_voter(41));                                                                           
                tmr_registers(1)(42)    <= not(local_tmr_voter(41));                                                                           
                tmr_registers(2)(42)    <= not(local_tmr_voter(41));                                                                           
 
                tmr_registers(0)(43)    <= not(local_tmr_voter(42));                                                                           
                tmr_registers(1)(43)    <= not(local_tmr_voter(42));                                                                           
                tmr_registers(2)(43)    <= not(local_tmr_voter(42));                                                                           
 
                tmr_registers(0)(44)    <= not(local_tmr_voter(43));                                                                           
                tmr_registers(1)(44)    <= not(local_tmr_voter(43));                                                                           
                tmr_registers(2)(44)    <= not(local_tmr_voter(43));                                                                           
 
                tmr_registers(0)(45)    <= not(local_tmr_voter(44));                                                                           
                tmr_registers(1)(45)    <= not(local_tmr_voter(44));                                                                           
                tmr_registers(2)(45)    <= not(local_tmr_voter(44));                                                                           
 
                tmr_registers(0)(46)    <= not(local_tmr_voter(45));                                                                           
                tmr_registers(1)(46)    <= not(local_tmr_voter(45));                                                                           
                tmr_registers(2)(46)    <= not(local_tmr_voter(45));                                                                           
 
                tmr_registers(0)(47)    <= not(local_tmr_voter(46));                                                                           
                tmr_registers(1)(47)    <= not(local_tmr_voter(46));                                                                           
                tmr_registers(2)(47)    <= not(local_tmr_voter(46));                                                                           
 
                tmr_registers(0)(48)    <= not(local_tmr_voter(47));                                                                           
                tmr_registers(1)(48)    <= not(local_tmr_voter(47));                                                                           
                tmr_registers(2)(48)    <= not(local_tmr_voter(47));                                                                           
 
                tmr_registers(0)(49)    <= not(local_tmr_voter(48));                                                                           
                tmr_registers(1)(49)    <= not(local_tmr_voter(48));                                                                           
                tmr_registers(2)(49)    <= not(local_tmr_voter(48));                                                                           
 
                tmr_registers(0)(50)    <= not(local_tmr_voter(49));                                                                           
                tmr_registers(1)(50)    <= not(local_tmr_voter(49));                                                                           
                tmr_registers(2)(50)    <= not(local_tmr_voter(49));                                                                           
 
                tmr_registers(0)(51)    <= not(local_tmr_voter(50));                                                                           
                tmr_registers(1)(51)    <= not(local_tmr_voter(50));                                                                           
                tmr_registers(2)(51)    <= not(local_tmr_voter(50));                                                                           
 
                tmr_registers(0)(52)    <= not(local_tmr_voter(51));                                                                           
                tmr_registers(1)(52)    <= not(local_tmr_voter(51));                                                                           
                tmr_registers(2)(52)    <= not(local_tmr_voter(51));                                                                           
 
                tmr_registers(0)(53)    <= not(local_tmr_voter(52));                                                                           
                tmr_registers(1)(53)    <= not(local_tmr_voter(52));                                                                           
                tmr_registers(2)(53)    <= not(local_tmr_voter(52));                                                                           
 
                tmr_registers(0)(54)    <= not(local_tmr_voter(53));                                                                           
                tmr_registers(1)(54)    <= not(local_tmr_voter(53));                                                                           
                tmr_registers(2)(54)    <= not(local_tmr_voter(53));                                                                           
 
                tmr_registers(0)(55)    <= not(local_tmr_voter(54));                                                                           
                tmr_registers(1)(55)    <= not(local_tmr_voter(54));                                                                           
                tmr_registers(2)(55)    <= not(local_tmr_voter(54));                                                                           
 
                tmr_registers(0)(56)    <= not(local_tmr_voter(55));                                                                           
                tmr_registers(1)(56)    <= not(local_tmr_voter(55));                                                                           
                tmr_registers(2)(56)    <= not(local_tmr_voter(55));                                                                           
 
                tmr_registers(0)(57)    <= not(local_tmr_voter(56));                                                                           
                tmr_registers(1)(57)    <= not(local_tmr_voter(56));                                                                           
                tmr_registers(2)(57)    <= not(local_tmr_voter(56));                                                                           
 
                tmr_registers(0)(58)    <= not(local_tmr_voter(57));                                                                           
                tmr_registers(1)(58)    <= not(local_tmr_voter(57));                                                                           
                tmr_registers(2)(58)    <= not(local_tmr_voter(57));                                                                           
 
                tmr_registers(0)(59)    <= not(local_tmr_voter(58));                                                                           
                tmr_registers(1)(59)    <= not(local_tmr_voter(58));                                                                           
                tmr_registers(2)(59)    <= not(local_tmr_voter(58));                                                                           
 
                tmr_registers(0)(60)    <= not(local_tmr_voter(59));                                                                           
                tmr_registers(1)(60)    <= not(local_tmr_voter(59));                                                                           
                tmr_registers(2)(60)    <= not(local_tmr_voter(59));                                                                           
 
                tmr_registers(0)(61)    <= not(local_tmr_voter(60));                                                                           
                tmr_registers(1)(61)    <= not(local_tmr_voter(60));                                                                           
                tmr_registers(2)(61)    <= not(local_tmr_voter(60));                                                                           
 
                tmr_registers(0)(62)    <= not(local_tmr_voter(61));                                                                           
                tmr_registers(1)(62)    <= not(local_tmr_voter(61));                                                                           
                tmr_registers(2)(62)    <= not(local_tmr_voter(61));                                                                           
 
                tmr_registers(0)(63)    <= not(local_tmr_voter(62));                                                                           
                tmr_registers(1)(63)    <= not(local_tmr_voter(62));                                                                           
                tmr_registers(2)(63)    <= not(local_tmr_voter(62));                                                                           
 
                tmr_registers(0)(64)    <= not(local_tmr_voter(63));                                                                           
                tmr_registers(1)(64)    <= not(local_tmr_voter(63));                                                                           
                tmr_registers(2)(64)    <= not(local_tmr_voter(63));                                                                           
 
                tmr_registers(0)(65)    <= not(local_tmr_voter(64));                                                                           
                tmr_registers(1)(65)    <= not(local_tmr_voter(64));                                                                           
                tmr_registers(2)(65)    <= not(local_tmr_voter(64));                                                                           
 
                tmr_registers(0)(66)    <= not(local_tmr_voter(65));                                                                           
                tmr_registers(1)(66)    <= not(local_tmr_voter(65));                                                                           
                tmr_registers(2)(66)    <= not(local_tmr_voter(65));                                                                           
 
                tmr_registers(0)(67)    <= not(local_tmr_voter(66));                                                                           
                tmr_registers(1)(67)    <= not(local_tmr_voter(66));                                                                           
                tmr_registers(2)(67)    <= not(local_tmr_voter(66));                                                                           
 
                tmr_registers(0)(68)    <= not(local_tmr_voter(67));                                                                           
                tmr_registers(1)(68)    <= not(local_tmr_voter(67));                                                                           
                tmr_registers(2)(68)    <= not(local_tmr_voter(67));                                                                           
 
                tmr_registers(0)(69)    <= not(local_tmr_voter(68));                                                                           
                tmr_registers(1)(69)    <= not(local_tmr_voter(68));                                                                           
                tmr_registers(2)(69)    <= not(local_tmr_voter(68));                                                                           
 
                tmr_registers(0)(70)    <= not(local_tmr_voter(69));                                                                           
                tmr_registers(1)(70)    <= not(local_tmr_voter(69));                                                                           
                tmr_registers(2)(70)    <= not(local_tmr_voter(69));                                                                           
 
                tmr_registers(0)(71)    <= not(local_tmr_voter(70));                                                                           
                tmr_registers(1)(71)    <= not(local_tmr_voter(70));                                                                           
                tmr_registers(2)(71)    <= not(local_tmr_voter(70));                                                                           
 
                tmr_registers(0)(72)    <= not(local_tmr_voter(71));                                                                           
                tmr_registers(1)(72)    <= not(local_tmr_voter(71));                                                                           
                tmr_registers(2)(72)    <= not(local_tmr_voter(71));                                                                           
 
                tmr_registers(0)(73)    <= not(local_tmr_voter(72));                                                                           
                tmr_registers(1)(73)    <= not(local_tmr_voter(72));                                                                           
                tmr_registers(2)(73)    <= not(local_tmr_voter(72));                                                                           
 
                tmr_registers(0)(74)    <= not(local_tmr_voter(73));                                                                           
                tmr_registers(1)(74)    <= not(local_tmr_voter(73));                                                                           
                tmr_registers(2)(74)    <= not(local_tmr_voter(73));                                                                           
 
                tmr_registers(0)(75)    <= not(local_tmr_voter(74));                                                                           
                tmr_registers(1)(75)    <= not(local_tmr_voter(74));                                                                           
                tmr_registers(2)(75)    <= not(local_tmr_voter(74));                                                                           
 
                tmr_registers(0)(76)    <= not(local_tmr_voter(75));                                                                           
                tmr_registers(1)(76)    <= not(local_tmr_voter(75));                                                                           
                tmr_registers(2)(76)    <= not(local_tmr_voter(75));                                                                           
 
                tmr_registers(0)(77)    <= not(local_tmr_voter(76));                                                                           
                tmr_registers(1)(77)    <= not(local_tmr_voter(76));                                                                           
                tmr_registers(2)(77)    <= not(local_tmr_voter(76));                                                                           
 
                tmr_registers(0)(78)    <= not(local_tmr_voter(77));                                                                           
                tmr_registers(1)(78)    <= not(local_tmr_voter(77));                                                                           
                tmr_registers(2)(78)    <= not(local_tmr_voter(77));                                                                           
 
                tmr_registers(0)(79)    <= not(local_tmr_voter(78));                                                                           
                tmr_registers(1)(79)    <= not(local_tmr_voter(78));                                                                           
                tmr_registers(2)(79)    <= not(local_tmr_voter(78));                                                                           
 
                tmr_registers(0)(80)    <= not(local_tmr_voter(79));                                                                           
                tmr_registers(1)(80)    <= not(local_tmr_voter(79));                                                                           
                tmr_registers(2)(80)    <= not(local_tmr_voter(79));                                                                           
 
                tmr_registers(0)(81)    <= not(local_tmr_voter(80));                                                                           
                tmr_registers(1)(81)    <= not(local_tmr_voter(80));                                                                           
                tmr_registers(2)(81)    <= not(local_tmr_voter(80));                                                                           
 
                tmr_registers(0)(82)    <= not(local_tmr_voter(81));                                                                           
                tmr_registers(1)(82)    <= not(local_tmr_voter(81));                                                                           
                tmr_registers(2)(82)    <= not(local_tmr_voter(81));                                                                           
 
                tmr_registers(0)(83)    <= not(local_tmr_voter(82));                                                                           
                tmr_registers(1)(83)    <= not(local_tmr_voter(82));                                                                           
                tmr_registers(2)(83)    <= not(local_tmr_voter(82));                                                                           
 
                tmr_registers(0)(84)    <= not(local_tmr_voter(83));                                                                           
                tmr_registers(1)(84)    <= not(local_tmr_voter(83));                                                                           
                tmr_registers(2)(84)    <= not(local_tmr_voter(83));                                                                           
 
                tmr_registers(0)(85)    <= not(local_tmr_voter(84));                                                                           
                tmr_registers(1)(85)    <= not(local_tmr_voter(84));                                                                           
                tmr_registers(2)(85)    <= not(local_tmr_voter(84));                                                                           
 
                tmr_registers(0)(86)    <= not(local_tmr_voter(85));                                                                           
                tmr_registers(1)(86)    <= not(local_tmr_voter(85));                                                                           
                tmr_registers(2)(86)    <= not(local_tmr_voter(85));                                                                           
 
                tmr_registers(0)(87)    <= not(local_tmr_voter(86));                                                                           
                tmr_registers(1)(87)    <= not(local_tmr_voter(86));                                                                           
                tmr_registers(2)(87)    <= not(local_tmr_voter(86));                                                                           
 
                tmr_registers(0)(88)    <= not(local_tmr_voter(87));                                                                           
                tmr_registers(1)(88)    <= not(local_tmr_voter(87));                                                                           
                tmr_registers(2)(88)    <= not(local_tmr_voter(87));                                                                           
 
                tmr_registers(0)(89)    <= not(local_tmr_voter(88));                                                                           
                tmr_registers(1)(89)    <= not(local_tmr_voter(88));                                                                           
                tmr_registers(2)(89)    <= not(local_tmr_voter(88));                                                                           
 
                tmr_registers(0)(90)    <= not(local_tmr_voter(89));                                                                           
                tmr_registers(1)(90)    <= not(local_tmr_voter(89));                                                                           
                tmr_registers(2)(90)    <= not(local_tmr_voter(89));                                                                           
 
                tmr_registers(0)(91)    <= not(local_tmr_voter(90));                                                                           
                tmr_registers(1)(91)    <= not(local_tmr_voter(90));                                                                           
                tmr_registers(2)(91)    <= not(local_tmr_voter(90));                                                                           
 
                tmr_registers(0)(92)    <= not(local_tmr_voter(91));                                                                           
                tmr_registers(1)(92)    <= not(local_tmr_voter(91));                                                                           
                tmr_registers(2)(92)    <= not(local_tmr_voter(91));                                                                           
 
                tmr_registers(0)(93)    <= not(local_tmr_voter(92));                                                                           
                tmr_registers(1)(93)    <= not(local_tmr_voter(92));                                                                           
                tmr_registers(2)(93)    <= not(local_tmr_voter(92));                                                                           
 
                tmr_registers(0)(94)    <= not(local_tmr_voter(93));                                                                           
                tmr_registers(1)(94)    <= not(local_tmr_voter(93));                                                                           
                tmr_registers(2)(94)    <= not(local_tmr_voter(93));                                                                           
 
                tmr_registers(0)(95)    <= not(local_tmr_voter(94));                                                                           
                tmr_registers(1)(95)    <= not(local_tmr_voter(94));                                                                           
                tmr_registers(2)(95)    <= not(local_tmr_voter(94));                                                                           
 
                tmr_registers(0)(96)    <= not(local_tmr_voter(95));                                                                           
                tmr_registers(1)(96)    <= not(local_tmr_voter(95));                                                                           
                tmr_registers(2)(96)    <= not(local_tmr_voter(95));                                                                           
 
                tmr_registers(0)(97)    <= not(local_tmr_voter(96));                                                                           
                tmr_registers(1)(97)    <= not(local_tmr_voter(96));                                                                           
                tmr_registers(2)(97)    <= not(local_tmr_voter(96));                                                                           
 
                tmr_registers(0)(98)    <= not(local_tmr_voter(97));                                                                           
                tmr_registers(1)(98)    <= not(local_tmr_voter(97));                                                                           
                tmr_registers(2)(98)    <= not(local_tmr_voter(97));                                                                           
 
                tmr_registers(0)(99)    <= not(local_tmr_voter(98));                                                                           
                tmr_registers(1)(99)    <= not(local_tmr_voter(98));                                                                           
                tmr_registers(2)(99)    <= not(local_tmr_voter(98));                                                                           
 
                tmr_registers(0)(100)    <= not(local_tmr_voter(99));                                                                           
                tmr_registers(1)(100)    <= not(local_tmr_voter(99));                                                                           
                tmr_registers(2)(100)    <= not(local_tmr_voter(99));                                                                           
 
                tmr_registers(0)(101)    <= not(local_tmr_voter(100));                                                                           
                tmr_registers(1)(101)    <= not(local_tmr_voter(100));                                                                           
                tmr_registers(2)(101)    <= not(local_tmr_voter(100));                                                                           
 
                tmr_registers(0)(102)    <= not(local_tmr_voter(101));                                                                           
                tmr_registers(1)(102)    <= not(local_tmr_voter(101));                                                                           
                tmr_registers(2)(102)    <= not(local_tmr_voter(101));                                                                           
 
                tmr_registers(0)(103)    <= not(local_tmr_voter(102));                                                                           
                tmr_registers(1)(103)    <= not(local_tmr_voter(102));                                                                           
                tmr_registers(2)(103)    <= not(local_tmr_voter(102));                                                                           
 
                tmr_registers(0)(104)    <= not(local_tmr_voter(103));                                                                           
                tmr_registers(1)(104)    <= not(local_tmr_voter(103));                                                                           
                tmr_registers(2)(104)    <= not(local_tmr_voter(103));                                                                           
 
                tmr_registers(0)(105)    <= not(local_tmr_voter(104));                                                                           
                tmr_registers(1)(105)    <= not(local_tmr_voter(104));                                                                           
                tmr_registers(2)(105)    <= not(local_tmr_voter(104));                                                                           
 
                tmr_registers(0)(106)    <= not(local_tmr_voter(105));                                                                           
                tmr_registers(1)(106)    <= not(local_tmr_voter(105));                                                                           
                tmr_registers(2)(106)    <= not(local_tmr_voter(105));                                                                           
 
                tmr_registers(0)(107)    <= not(local_tmr_voter(106));                                                                           
                tmr_registers(1)(107)    <= not(local_tmr_voter(106));                                                                           
                tmr_registers(2)(107)    <= not(local_tmr_voter(106));                                                                           
 
                tmr_registers(0)(108)    <= not(local_tmr_voter(107));                                                                           
                tmr_registers(1)(108)    <= not(local_tmr_voter(107));                                                                           
                tmr_registers(2)(108)    <= not(local_tmr_voter(107));                                                                           
 
                tmr_registers(0)(109)    <= not(local_tmr_voter(108));                                                                           
                tmr_registers(1)(109)    <= not(local_tmr_voter(108));                                                                           
                tmr_registers(2)(109)    <= not(local_tmr_voter(108));                                                                           
 
                tmr_registers(0)(110)    <= not(local_tmr_voter(109));                                                                           
                tmr_registers(1)(110)    <= not(local_tmr_voter(109));                                                                           
                tmr_registers(2)(110)    <= not(local_tmr_voter(109));                                                                           
 
                tmr_registers(0)(111)    <= not(local_tmr_voter(110));                                                                           
                tmr_registers(1)(111)    <= not(local_tmr_voter(110));                                                                           
                tmr_registers(2)(111)    <= not(local_tmr_voter(110));                                                                           
 
                tmr_registers(0)(112)    <= not(local_tmr_voter(111));                                                                           
                tmr_registers(1)(112)    <= not(local_tmr_voter(111));                                                                           
                tmr_registers(2)(112)    <= not(local_tmr_voter(111));                                                                           
 
                tmr_registers(0)(113)    <= not(local_tmr_voter(112));                                                                           
                tmr_registers(1)(113)    <= not(local_tmr_voter(112));                                                                           
                tmr_registers(2)(113)    <= not(local_tmr_voter(112));                                                                           
 
                tmr_registers(0)(114)    <= not(local_tmr_voter(113));                                                                           
                tmr_registers(1)(114)    <= not(local_tmr_voter(113));                                                                           
                tmr_registers(2)(114)    <= not(local_tmr_voter(113));                                                                           
 
                tmr_registers(0)(115)    <= not(local_tmr_voter(114));                                                                           
                tmr_registers(1)(115)    <= not(local_tmr_voter(114));                                                                           
                tmr_registers(2)(115)    <= not(local_tmr_voter(114));                                                                           
 
                tmr_registers(0)(116)    <= not(local_tmr_voter(115));                                                                           
                tmr_registers(1)(116)    <= not(local_tmr_voter(115));                                                                           
                tmr_registers(2)(116)    <= not(local_tmr_voter(115));                                                                           
 
                tmr_registers(0)(117)    <= not(local_tmr_voter(116));                                                                           
                tmr_registers(1)(117)    <= not(local_tmr_voter(116));                                                                           
                tmr_registers(2)(117)    <= not(local_tmr_voter(116));                                                                           
 
                tmr_registers(0)(118)    <= not(local_tmr_voter(117));                                                                           
                tmr_registers(1)(118)    <= not(local_tmr_voter(117));                                                                           
                tmr_registers(2)(118)    <= not(local_tmr_voter(117));                                                                           
 
                tmr_registers(0)(119)    <= not(local_tmr_voter(118));                                                                           
                tmr_registers(1)(119)    <= not(local_tmr_voter(118));                                                                           
                tmr_registers(2)(119)    <= not(local_tmr_voter(118));                                                                           
 
                tmr_registers(0)(120)    <= not(local_tmr_voter(119));                                                                           
                tmr_registers(1)(120)    <= not(local_tmr_voter(119));                                                                           
                tmr_registers(2)(120)    <= not(local_tmr_voter(119));                                                                           
 
                tmr_registers(0)(121)    <= not(local_tmr_voter(120));                                                                           
                tmr_registers(1)(121)    <= not(local_tmr_voter(120));                                                                           
                tmr_registers(2)(121)    <= not(local_tmr_voter(120));                                                                           
 
                tmr_registers(0)(122)    <= not(local_tmr_voter(121));                                                                           
                tmr_registers(1)(122)    <= not(local_tmr_voter(121));                                                                           
                tmr_registers(2)(122)    <= not(local_tmr_voter(121));                                                                           
 
                tmr_registers(0)(123)    <= not(local_tmr_voter(122));                                                                           
                tmr_registers(1)(123)    <= not(local_tmr_voter(122));                                                                           
                tmr_registers(2)(123)    <= not(local_tmr_voter(122));                                                                           
 
                tmr_registers(0)(124)    <= not(local_tmr_voter(123));                                                                           
                tmr_registers(1)(124)    <= not(local_tmr_voter(123));                                                                           
                tmr_registers(2)(124)    <= not(local_tmr_voter(123));                                                                           
 
                tmr_registers(0)(125)    <= not(local_tmr_voter(124));                                                                           
                tmr_registers(1)(125)    <= not(local_tmr_voter(124));                                                                           
                tmr_registers(2)(125)    <= not(local_tmr_voter(124));                                                                           
 
                tmr_registers(0)(126)    <= not(local_tmr_voter(125));                                                                           
                tmr_registers(1)(126)    <= not(local_tmr_voter(125));                                                                           
                tmr_registers(2)(126)    <= not(local_tmr_voter(125));                                                                           
 
                tmr_registers(0)(127)    <= not(local_tmr_voter(126));                                                                           
                tmr_registers(1)(127)    <= not(local_tmr_voter(126));                                                                           
                tmr_registers(2)(127)    <= not(local_tmr_voter(126));                                                                           
 
                tmr_registers(0)(128)    <= not(local_tmr_voter(127));                                                                           
                tmr_registers(1)(128)    <= not(local_tmr_voter(127));                                                                           
                tmr_registers(2)(128)    <= not(local_tmr_voter(127));                                                                           
 
                tmr_registers(0)(129)    <= not(local_tmr_voter(128));                                                                           
                tmr_registers(1)(129)    <= not(local_tmr_voter(128));                                                                           
                tmr_registers(2)(129)    <= not(local_tmr_voter(128));                                                                           
 
                tmr_registers(0)(130)    <= not(local_tmr_voter(129));                                                                           
                tmr_registers(1)(130)    <= not(local_tmr_voter(129));                                                                           
                tmr_registers(2)(130)    <= not(local_tmr_voter(129));                                                                           
 
                tmr_registers(0)(131)    <= not(local_tmr_voter(130));                                                                           
                tmr_registers(1)(131)    <= not(local_tmr_voter(130));                                                                           
                tmr_registers(2)(131)    <= not(local_tmr_voter(130));                                                                           
 
                tmr_registers(0)(132)    <= not(local_tmr_voter(131));                                                                           
                tmr_registers(1)(132)    <= not(local_tmr_voter(131));                                                                           
                tmr_registers(2)(132)    <= not(local_tmr_voter(131));                                                                           
 
                tmr_registers(0)(133)    <= not(local_tmr_voter(132));                                                                           
                tmr_registers(1)(133)    <= not(local_tmr_voter(132));                                                                           
                tmr_registers(2)(133)    <= not(local_tmr_voter(132));                                                                           
 
                tmr_registers(0)(134)    <= not(local_tmr_voter(133));                                                                           
                tmr_registers(1)(134)    <= not(local_tmr_voter(133));                                                                           
                tmr_registers(2)(134)    <= not(local_tmr_voter(133));                                                                           
 
                tmr_registers(0)(135)    <= not(local_tmr_voter(134));                                                                           
                tmr_registers(1)(135)    <= not(local_tmr_voter(134));                                                                           
                tmr_registers(2)(135)    <= not(local_tmr_voter(134));                                                                           
 
                tmr_registers(0)(136)    <= not(local_tmr_voter(135));                                                                           
                tmr_registers(1)(136)    <= not(local_tmr_voter(135));                                                                           
                tmr_registers(2)(136)    <= not(local_tmr_voter(135));                                                                           
 
                tmr_registers(0)(137)    <= not(local_tmr_voter(136));                                                                           
                tmr_registers(1)(137)    <= not(local_tmr_voter(136));                                                                           
                tmr_registers(2)(137)    <= not(local_tmr_voter(136));                                                                           
 
                tmr_registers(0)(138)    <= not(local_tmr_voter(137));                                                                           
                tmr_registers(1)(138)    <= not(local_tmr_voter(137));                                                                           
                tmr_registers(2)(138)    <= not(local_tmr_voter(137));                                                                           
 
                tmr_registers(0)(139)    <= not(local_tmr_voter(138));                                                                           
                tmr_registers(1)(139)    <= not(local_tmr_voter(138));                                                                           
                tmr_registers(2)(139)    <= not(local_tmr_voter(138));                                                                           
 
                tmr_registers(0)(140)    <= not(local_tmr_voter(139));                                                                           
                tmr_registers(1)(140)    <= not(local_tmr_voter(139));                                                                           
                tmr_registers(2)(140)    <= not(local_tmr_voter(139));                                                                           
 
                tmr_registers(0)(141)    <= not(local_tmr_voter(140));                                                                           
                tmr_registers(1)(141)    <= not(local_tmr_voter(140));                                                                           
                tmr_registers(2)(141)    <= not(local_tmr_voter(140));                                                                           
 
                tmr_registers(0)(142)    <= not(local_tmr_voter(141));                                                                           
                tmr_registers(1)(142)    <= not(local_tmr_voter(141));                                                                           
                tmr_registers(2)(142)    <= not(local_tmr_voter(141));                                                                           
 
                tmr_registers(0)(143)    <= not(local_tmr_voter(142));                                                                           
                tmr_registers(1)(143)    <= not(local_tmr_voter(142));                                                                           
                tmr_registers(2)(143)    <= not(local_tmr_voter(142));                                                                           
 
                tmr_registers(0)(144)    <= not(local_tmr_voter(143));                                                                           
                tmr_registers(1)(144)    <= not(local_tmr_voter(143));                                                                           
                tmr_registers(2)(144)    <= not(local_tmr_voter(143));                                                                           
 
                tmr_registers(0)(145)    <= not(local_tmr_voter(144));                                                                           
                tmr_registers(1)(145)    <= not(local_tmr_voter(144));                                                                           
                tmr_registers(2)(145)    <= not(local_tmr_voter(144));                                                                           
 
                tmr_registers(0)(146)    <= not(local_tmr_voter(145));                                                                           
                tmr_registers(1)(146)    <= not(local_tmr_voter(145));                                                                           
                tmr_registers(2)(146)    <= not(local_tmr_voter(145));                                                                           
 
                tmr_registers(0)(147)    <= not(local_tmr_voter(146));                                                                           
                tmr_registers(1)(147)    <= not(local_tmr_voter(146));                                                                           
                tmr_registers(2)(147)    <= not(local_tmr_voter(146));                                                                           
 
                tmr_registers(0)(148)    <= not(local_tmr_voter(147));                                                                           
                tmr_registers(1)(148)    <= not(local_tmr_voter(147));                                                                           
                tmr_registers(2)(148)    <= not(local_tmr_voter(147));                                                                           
 
                tmr_registers(0)(149)    <= not(local_tmr_voter(148));                                                                           
                tmr_registers(1)(149)    <= not(local_tmr_voter(148));                                                                           
                tmr_registers(2)(149)    <= not(local_tmr_voter(148));                                                                           
 
                tmr_registers(0)(150)    <= not(local_tmr_voter(149));                                                                           
                tmr_registers(1)(150)    <= not(local_tmr_voter(149));                                                                           
                tmr_registers(2)(150)    <= not(local_tmr_voter(149));                                                                           
 
                tmr_registers(0)(151)    <= not(local_tmr_voter(150));                                                                           
                tmr_registers(1)(151)    <= not(local_tmr_voter(150));                                                                           
                tmr_registers(2)(151)    <= not(local_tmr_voter(150));                                                                           
 
                tmr_registers(0)(152)    <= not(local_tmr_voter(151));                                                                           
                tmr_registers(1)(152)    <= not(local_tmr_voter(151));                                                                           
                tmr_registers(2)(152)    <= not(local_tmr_voter(151));                                                                           
 
                tmr_registers(0)(153)    <= not(local_tmr_voter(152));                                                                           
                tmr_registers(1)(153)    <= not(local_tmr_voter(152));                                                                           
                tmr_registers(2)(153)    <= not(local_tmr_voter(152));                                                                           
 
                tmr_registers(0)(154)    <= not(local_tmr_voter(153));                                                                           
                tmr_registers(1)(154)    <= not(local_tmr_voter(153));                                                                           
                tmr_registers(2)(154)    <= not(local_tmr_voter(153));                                                                           
 
                tmr_registers(0)(155)    <= not(local_tmr_voter(154));                                                                           
                tmr_registers(1)(155)    <= not(local_tmr_voter(154));                                                                           
                tmr_registers(2)(155)    <= not(local_tmr_voter(154));                                                                           
 
                tmr_registers(0)(156)    <= not(local_tmr_voter(155));                                                                           
                tmr_registers(1)(156)    <= not(local_tmr_voter(155));                                                                           
                tmr_registers(2)(156)    <= not(local_tmr_voter(155));                                                                           
 
                tmr_registers(0)(157)    <= not(local_tmr_voter(156));                                                                           
                tmr_registers(1)(157)    <= not(local_tmr_voter(156));                                                                           
                tmr_registers(2)(157)    <= not(local_tmr_voter(156));                                                                           
 
                tmr_registers(0)(158)    <= not(local_tmr_voter(157));                                                                           
                tmr_registers(1)(158)    <= not(local_tmr_voter(157));                                                                           
                tmr_registers(2)(158)    <= not(local_tmr_voter(157));                                                                           
 
                tmr_registers(0)(159)    <= not(local_tmr_voter(158));                                                                           
                tmr_registers(1)(159)    <= not(local_tmr_voter(158));                                                                           
                tmr_registers(2)(159)    <= not(local_tmr_voter(158));                                                                           
 
                tmr_registers(0)(160)    <= not(local_tmr_voter(159));                                                                           
                tmr_registers(1)(160)    <= not(local_tmr_voter(159));                                                                           
                tmr_registers(2)(160)    <= not(local_tmr_voter(159));                                                                           
 
                tmr_registers(0)(161)    <= not(local_tmr_voter(160));                                                                           
                tmr_registers(1)(161)    <= not(local_tmr_voter(160));                                                                           
                tmr_registers(2)(161)    <= not(local_tmr_voter(160));                                                                           
 
                tmr_registers(0)(162)    <= not(local_tmr_voter(161));                                                                           
                tmr_registers(1)(162)    <= not(local_tmr_voter(161));                                                                           
                tmr_registers(2)(162)    <= not(local_tmr_voter(161));                                                                           
 
                tmr_registers(0)(163)    <= not(local_tmr_voter(162));                                                                           
                tmr_registers(1)(163)    <= not(local_tmr_voter(162));                                                                           
                tmr_registers(2)(163)    <= not(local_tmr_voter(162));                                                                           
 
                tmr_registers(0)(164)    <= not(local_tmr_voter(163));                                                                           
                tmr_registers(1)(164)    <= not(local_tmr_voter(163));                                                                           
                tmr_registers(2)(164)    <= not(local_tmr_voter(163));                                                                           
 
                tmr_registers(0)(165)    <= not(local_tmr_voter(164));                                                                           
                tmr_registers(1)(165)    <= not(local_tmr_voter(164));                                                                           
                tmr_registers(2)(165)    <= not(local_tmr_voter(164));                                                                           
 
                tmr_registers(0)(166)    <= not(local_tmr_voter(165));                                                                           
                tmr_registers(1)(166)    <= not(local_tmr_voter(165));                                                                           
                tmr_registers(2)(166)    <= not(local_tmr_voter(165));                                                                           
 
                tmr_registers(0)(167)    <= not(local_tmr_voter(166));                                                                           
                tmr_registers(1)(167)    <= not(local_tmr_voter(166));                                                                           
                tmr_registers(2)(167)    <= not(local_tmr_voter(166));                                                                           
 
                tmr_registers(0)(168)    <= not(local_tmr_voter(167));                                                                           
                tmr_registers(1)(168)    <= not(local_tmr_voter(167));                                                                           
                tmr_registers(2)(168)    <= not(local_tmr_voter(167));                                                                           
 
                tmr_registers(0)(169)    <= not(local_tmr_voter(168));                                                                           
                tmr_registers(1)(169)    <= not(local_tmr_voter(168));                                                                           
                tmr_registers(2)(169)    <= not(local_tmr_voter(168));                                                                           
 
                tmr_registers(0)(170)    <= not(local_tmr_voter(169));                                                                           
                tmr_registers(1)(170)    <= not(local_tmr_voter(169));                                                                           
                tmr_registers(2)(170)    <= not(local_tmr_voter(169));                                                                           
 
                tmr_registers(0)(171)    <= not(local_tmr_voter(170));                                                                           
                tmr_registers(1)(171)    <= not(local_tmr_voter(170));                                                                           
                tmr_registers(2)(171)    <= not(local_tmr_voter(170));                                                                           
 
                tmr_registers(0)(172)    <= not(local_tmr_voter(171));                                                                           
                tmr_registers(1)(172)    <= not(local_tmr_voter(171));                                                                           
                tmr_registers(2)(172)    <= not(local_tmr_voter(171));                                                                           
 
                tmr_registers(0)(173)    <= not(local_tmr_voter(172));                                                                           
                tmr_registers(1)(173)    <= not(local_tmr_voter(172));                                                                           
                tmr_registers(2)(173)    <= not(local_tmr_voter(172));                                                                           
 
                tmr_registers(0)(174)    <= not(local_tmr_voter(173));                                                                           
                tmr_registers(1)(174)    <= not(local_tmr_voter(173));                                                                           
                tmr_registers(2)(174)    <= not(local_tmr_voter(173));                                                                           
 
                tmr_registers(0)(175)    <= not(local_tmr_voter(174));                                                                           
                tmr_registers(1)(175)    <= not(local_tmr_voter(174));                                                                           
                tmr_registers(2)(175)    <= not(local_tmr_voter(174));                                                                           
 
                tmr_registers(0)(176)    <= not(local_tmr_voter(175));                                                                           
                tmr_registers(1)(176)    <= not(local_tmr_voter(175));                                                                           
                tmr_registers(2)(176)    <= not(local_tmr_voter(175));                                                                           
 
                tmr_registers(0)(177)    <= not(local_tmr_voter(176));                                                                           
                tmr_registers(1)(177)    <= not(local_tmr_voter(176));                                                                           
                tmr_registers(2)(177)    <= not(local_tmr_voter(176));                                                                           
 
                tmr_registers(0)(178)    <= not(local_tmr_voter(177));                                                                           
                tmr_registers(1)(178)    <= not(local_tmr_voter(177));                                                                           
                tmr_registers(2)(178)    <= not(local_tmr_voter(177));                                                                           
 
                tmr_registers(0)(179)    <= not(local_tmr_voter(178));                                                                           
                tmr_registers(1)(179)    <= not(local_tmr_voter(178));                                                                           
                tmr_registers(2)(179)    <= not(local_tmr_voter(178));                                                                           
 
                tmr_registers(0)(180)    <= not(local_tmr_voter(179));                                                                           
                tmr_registers(1)(180)    <= not(local_tmr_voter(179));                                                                           
                tmr_registers(2)(180)    <= not(local_tmr_voter(179));                                                                           
 
                tmr_registers(0)(181)    <= not(local_tmr_voter(180));                                                                           
                tmr_registers(1)(181)    <= not(local_tmr_voter(180));                                                                           
                tmr_registers(2)(181)    <= not(local_tmr_voter(180));                                                                           
 
                tmr_registers(0)(182)    <= not(local_tmr_voter(181));                                                                           
                tmr_registers(1)(182)    <= not(local_tmr_voter(181));                                                                           
                tmr_registers(2)(182)    <= not(local_tmr_voter(181));                                                                           
 
                tmr_registers(0)(183)    <= not(local_tmr_voter(182));                                                                           
                tmr_registers(1)(183)    <= not(local_tmr_voter(182));                                                                           
                tmr_registers(2)(183)    <= not(local_tmr_voter(182));                                                                           
 
                tmr_registers(0)(184)    <= not(local_tmr_voter(183));                                                                           
                tmr_registers(1)(184)    <= not(local_tmr_voter(183));                                                                           
                tmr_registers(2)(184)    <= not(local_tmr_voter(183));                                                                           
 
                tmr_registers(0)(185)    <= not(local_tmr_voter(184));                                                                           
                tmr_registers(1)(185)    <= not(local_tmr_voter(184));                                                                           
                tmr_registers(2)(185)    <= not(local_tmr_voter(184));                                                                           
 
                tmr_registers(0)(186)    <= not(local_tmr_voter(185));                                                                           
                tmr_registers(1)(186)    <= not(local_tmr_voter(185));                                                                           
                tmr_registers(2)(186)    <= not(local_tmr_voter(185));                                                                           
 
                tmr_registers(0)(187)    <= not(local_tmr_voter(186));                                                                           
                tmr_registers(1)(187)    <= not(local_tmr_voter(186));                                                                           
                tmr_registers(2)(187)    <= not(local_tmr_voter(186));                                                                           
 
                tmr_registers(0)(188)    <= not(local_tmr_voter(187));                                                                           
                tmr_registers(1)(188)    <= not(local_tmr_voter(187));                                                                           
                tmr_registers(2)(188)    <= not(local_tmr_voter(187));                                                                           
 
                tmr_registers(0)(189)    <= not(local_tmr_voter(188));                                                                           
                tmr_registers(1)(189)    <= not(local_tmr_voter(188));                                                                           
                tmr_registers(2)(189)    <= not(local_tmr_voter(188));                                                                           
 
                tmr_registers(0)(190)    <= not(local_tmr_voter(189));                                                                           
                tmr_registers(1)(190)    <= not(local_tmr_voter(189));                                                                           
                tmr_registers(2)(190)    <= not(local_tmr_voter(189));                                                                           
 
                tmr_registers(0)(191)    <= not(local_tmr_voter(190));                                                                           
                tmr_registers(1)(191)    <= not(local_tmr_voter(190));                                                                           
                tmr_registers(2)(191)    <= not(local_tmr_voter(190));                                                                           
 
                tmr_registers(0)(192)    <= not(local_tmr_voter(191));                                                                           
                tmr_registers(1)(192)    <= not(local_tmr_voter(191));                                                                           
                tmr_registers(2)(192)    <= not(local_tmr_voter(191));                                                                           
 
                tmr_registers(0)(193)    <= not(local_tmr_voter(192));                                                                           
                tmr_registers(1)(193)    <= not(local_tmr_voter(192));                                                                           
                tmr_registers(2)(193)    <= not(local_tmr_voter(192));                                                                           
 
                tmr_registers(0)(194)    <= not(local_tmr_voter(193));                                                                           
                tmr_registers(1)(194)    <= not(local_tmr_voter(193));                                                                           
                tmr_registers(2)(194)    <= not(local_tmr_voter(193));                                                                           
 
                tmr_registers(0)(195)    <= not(local_tmr_voter(194));                                                                           
                tmr_registers(1)(195)    <= not(local_tmr_voter(194));                                                                           
                tmr_registers(2)(195)    <= not(local_tmr_voter(194));                                                                           
 
                tmr_registers(0)(196)    <= not(local_tmr_voter(195));                                                                           
                tmr_registers(1)(196)    <= not(local_tmr_voter(195));                                                                           
                tmr_registers(2)(196)    <= not(local_tmr_voter(195));                                                                           
 
                tmr_registers(0)(197)    <= not(local_tmr_voter(196));                                                                           
                tmr_registers(1)(197)    <= not(local_tmr_voter(196));                                                                           
                tmr_registers(2)(197)    <= not(local_tmr_voter(196));                                                                           
 
                tmr_registers(0)(198)    <= not(local_tmr_voter(197));                                                                           
                tmr_registers(1)(198)    <= not(local_tmr_voter(197));                                                                           
                tmr_registers(2)(198)    <= not(local_tmr_voter(197));                                                                           
 
                tmr_registers(0)(199)    <= not(local_tmr_voter(198));                                                                           
                tmr_registers(1)(199)    <= not(local_tmr_voter(198));                                                                           
                tmr_registers(2)(199)    <= not(local_tmr_voter(198));                                                                           
 
                tmr_registers(0)(200)    <= not(local_tmr_voter(199));                                                                           
                tmr_registers(1)(200)    <= not(local_tmr_voter(199));                                                                           
                tmr_registers(2)(200)    <= not(local_tmr_voter(199));                                                                           
 
                tmr_registers(0)(201)    <= not(local_tmr_voter(200));                                                                           
                tmr_registers(1)(201)    <= not(local_tmr_voter(200));                                                                           
                tmr_registers(2)(201)    <= not(local_tmr_voter(200));                                                                           
 
                tmr_registers(0)(202)    <= not(local_tmr_voter(201));                                                                           
                tmr_registers(1)(202)    <= not(local_tmr_voter(201));                                                                           
                tmr_registers(2)(202)    <= not(local_tmr_voter(201));                                                                           
 
                tmr_registers(0)(203)    <= not(local_tmr_voter(202));                                                                           
                tmr_registers(1)(203)    <= not(local_tmr_voter(202));                                                                           
                tmr_registers(2)(203)    <= not(local_tmr_voter(202));                                                                           
 
                tmr_registers(0)(204)    <= not(local_tmr_voter(203));                                                                           
                tmr_registers(1)(204)    <= not(local_tmr_voter(203));                                                                           
                tmr_registers(2)(204)    <= not(local_tmr_voter(203));                                                                           
 
                tmr_registers(0)(205)    <= not(local_tmr_voter(204));                                                                           
                tmr_registers(1)(205)    <= not(local_tmr_voter(204));                                                                           
                tmr_registers(2)(205)    <= not(local_tmr_voter(204));                                                                           
 
                tmr_registers(0)(206)    <= not(local_tmr_voter(205));                                                                           
                tmr_registers(1)(206)    <= not(local_tmr_voter(205));                                                                           
                tmr_registers(2)(206)    <= not(local_tmr_voter(205));                                                                           
 
                tmr_registers(0)(207)    <= not(local_tmr_voter(206));                                                                           
                tmr_registers(1)(207)    <= not(local_tmr_voter(206));                                                                           
                tmr_registers(2)(207)    <= not(local_tmr_voter(206));                                                                           
 
                tmr_registers(0)(208)    <= not(local_tmr_voter(207));                                                                           
                tmr_registers(1)(208)    <= not(local_tmr_voter(207));                                                                           
                tmr_registers(2)(208)    <= not(local_tmr_voter(207));                                                                           
 
                tmr_registers(0)(209)    <= not(local_tmr_voter(208));                                                                           
                tmr_registers(1)(209)    <= not(local_tmr_voter(208));                                                                           
                tmr_registers(2)(209)    <= not(local_tmr_voter(208));                                                                           
 
                tmr_registers(0)(210)    <= not(local_tmr_voter(209));                                                                           
                tmr_registers(1)(210)    <= not(local_tmr_voter(209));                                                                           
                tmr_registers(2)(210)    <= not(local_tmr_voter(209));                                                                           
 
                tmr_registers(0)(211)    <= not(local_tmr_voter(210));                                                                           
                tmr_registers(1)(211)    <= not(local_tmr_voter(210));                                                                           
                tmr_registers(2)(211)    <= not(local_tmr_voter(210));                                                                           
 
                tmr_registers(0)(212)    <= not(local_tmr_voter(211));                                                                           
                tmr_registers(1)(212)    <= not(local_tmr_voter(211));                                                                           
                tmr_registers(2)(212)    <= not(local_tmr_voter(211));                                                                           
 
                tmr_registers(0)(213)    <= not(local_tmr_voter(212));                                                                           
                tmr_registers(1)(213)    <= not(local_tmr_voter(212));                                                                           
                tmr_registers(2)(213)    <= not(local_tmr_voter(212));                                                                           
 
                tmr_registers(0)(214)    <= not(local_tmr_voter(213));                                                                           
                tmr_registers(1)(214)    <= not(local_tmr_voter(213));                                                                           
                tmr_registers(2)(214)    <= not(local_tmr_voter(213));                                                                           
 
                tmr_registers(0)(215)    <= not(local_tmr_voter(214));                                                                           
                tmr_registers(1)(215)    <= not(local_tmr_voter(214));                                                                           
                tmr_registers(2)(215)    <= not(local_tmr_voter(214));                                                                           
 
                tmr_registers(0)(216)    <= not(local_tmr_voter(215));                                                                           
                tmr_registers(1)(216)    <= not(local_tmr_voter(215));                                                                           
                tmr_registers(2)(216)    <= not(local_tmr_voter(215));                                                                           
 
                tmr_registers(0)(217)    <= not(local_tmr_voter(216));                                                                           
                tmr_registers(1)(217)    <= not(local_tmr_voter(216));                                                                           
                tmr_registers(2)(217)    <= not(local_tmr_voter(216));                                                                           
 
                tmr_registers(0)(218)    <= not(local_tmr_voter(217));                                                                           
                tmr_registers(1)(218)    <= not(local_tmr_voter(217));                                                                           
                tmr_registers(2)(218)    <= not(local_tmr_voter(217));                                                                           
 
                tmr_registers(0)(219)    <= not(local_tmr_voter(218));                                                                           
                tmr_registers(1)(219)    <= not(local_tmr_voter(218));                                                                           
                tmr_registers(2)(219)    <= not(local_tmr_voter(218));                                                                           
 
                tmr_registers(0)(220)    <= not(local_tmr_voter(219));                                                                           
                tmr_registers(1)(220)    <= not(local_tmr_voter(219));                                                                           
                tmr_registers(2)(220)    <= not(local_tmr_voter(219));                                                                           
 
                tmr_registers(0)(221)    <= not(local_tmr_voter(220));                                                                           
                tmr_registers(1)(221)    <= not(local_tmr_voter(220));                                                                           
                tmr_registers(2)(221)    <= not(local_tmr_voter(220));                                                                           
 
                tmr_registers(0)(222)    <= not(local_tmr_voter(221));                                                                           
                tmr_registers(1)(222)    <= not(local_tmr_voter(221));                                                                           
                tmr_registers(2)(222)    <= not(local_tmr_voter(221));                                                                           
 
                tmr_registers(0)(223)    <= not(local_tmr_voter(222));                                                                           
                tmr_registers(1)(223)    <= not(local_tmr_voter(222));                                                                           
                tmr_registers(2)(223)    <= not(local_tmr_voter(222));                                                                           
 
                tmr_registers(0)(224)    <= not(local_tmr_voter(223));                                                                           
                tmr_registers(1)(224)    <= not(local_tmr_voter(223));                                                                           
                tmr_registers(2)(224)    <= not(local_tmr_voter(223));                                                                           
 
                tmr_registers(0)(225)    <= not(local_tmr_voter(224));                                                                           
                tmr_registers(1)(225)    <= not(local_tmr_voter(224));                                                                           
                tmr_registers(2)(225)    <= not(local_tmr_voter(224));                                                                           
 
                tmr_registers(0)(226)    <= not(local_tmr_voter(225));                                                                           
                tmr_registers(1)(226)    <= not(local_tmr_voter(225));                                                                           
                tmr_registers(2)(226)    <= not(local_tmr_voter(225));                                                                           
 
                tmr_registers(0)(227)    <= not(local_tmr_voter(226));                                                                           
                tmr_registers(1)(227)    <= not(local_tmr_voter(226));                                                                           
                tmr_registers(2)(227)    <= not(local_tmr_voter(226));                                                                           
 
                tmr_registers(0)(228)    <= not(local_tmr_voter(227));                                                                           
                tmr_registers(1)(228)    <= not(local_tmr_voter(227));                                                                           
                tmr_registers(2)(228)    <= not(local_tmr_voter(227));                                                                           
 
                tmr_registers(0)(229)    <= not(local_tmr_voter(228));                                                                           
                tmr_registers(1)(229)    <= not(local_tmr_voter(228));                                                                           
                tmr_registers(2)(229)    <= not(local_tmr_voter(228));                                                                           
 
                tmr_registers(0)(230)    <= not(local_tmr_voter(229));                                                                           
                tmr_registers(1)(230)    <= not(local_tmr_voter(229));                                                                           
                tmr_registers(2)(230)    <= not(local_tmr_voter(229));                                                                           
 
                tmr_registers(0)(231)    <= not(local_tmr_voter(230));                                                                           
                tmr_registers(1)(231)    <= not(local_tmr_voter(230));                                                                           
                tmr_registers(2)(231)    <= not(local_tmr_voter(230));                                                                           
 
                tmr_registers(0)(232)    <= not(local_tmr_voter(231));                                                                           
                tmr_registers(1)(232)    <= not(local_tmr_voter(231));                                                                           
                tmr_registers(2)(232)    <= not(local_tmr_voter(231));                                                                           
 
                tmr_registers(0)(233)    <= not(local_tmr_voter(232));                                                                           
                tmr_registers(1)(233)    <= not(local_tmr_voter(232));                                                                           
                tmr_registers(2)(233)    <= not(local_tmr_voter(232));                                                                           
 
                tmr_registers(0)(234)    <= not(local_tmr_voter(233));                                                                           
                tmr_registers(1)(234)    <= not(local_tmr_voter(233));                                                                           
                tmr_registers(2)(234)    <= not(local_tmr_voter(233));                                                                           
 
                tmr_registers(0)(235)    <= not(local_tmr_voter(234));                                                                           
                tmr_registers(1)(235)    <= not(local_tmr_voter(234));                                                                           
                tmr_registers(2)(235)    <= not(local_tmr_voter(234));                                                                           
 
                tmr_registers(0)(236)    <= not(local_tmr_voter(235));                                                                           
                tmr_registers(1)(236)    <= not(local_tmr_voter(235));                                                                           
                tmr_registers(2)(236)    <= not(local_tmr_voter(235));                                                                           
 
                tmr_registers(0)(237)    <= not(local_tmr_voter(236));                                                                           
                tmr_registers(1)(237)    <= not(local_tmr_voter(236));                                                                           
                tmr_registers(2)(237)    <= not(local_tmr_voter(236));                                                                           
 
                tmr_registers(0)(238)    <= not(local_tmr_voter(237));                                                                           
                tmr_registers(1)(238)    <= not(local_tmr_voter(237));                                                                           
                tmr_registers(2)(238)    <= not(local_tmr_voter(237));                                                                           
 
                tmr_registers(0)(239)    <= not(local_tmr_voter(238));                                                                           
                tmr_registers(1)(239)    <= not(local_tmr_voter(238));                                                                           
                tmr_registers(2)(239)    <= not(local_tmr_voter(238));                                                                           
 
                tmr_registers(0)(240)    <= not(local_tmr_voter(239));                                                                           
                tmr_registers(1)(240)    <= not(local_tmr_voter(239));                                                                           
                tmr_registers(2)(240)    <= not(local_tmr_voter(239));                                                                           
 
                tmr_registers(0)(241)    <= not(local_tmr_voter(240));                                                                           
                tmr_registers(1)(241)    <= not(local_tmr_voter(240));                                                                           
                tmr_registers(2)(241)    <= not(local_tmr_voter(240));                                                                           
 
                tmr_registers(0)(242)    <= not(local_tmr_voter(241));                                                                           
                tmr_registers(1)(242)    <= not(local_tmr_voter(241));                                                                           
                tmr_registers(2)(242)    <= not(local_tmr_voter(241));                                                                           
 
                tmr_registers(0)(243)    <= not(local_tmr_voter(242));                                                                           
                tmr_registers(1)(243)    <= not(local_tmr_voter(242));                                                                           
                tmr_registers(2)(243)    <= not(local_tmr_voter(242));                                                                           
 
                tmr_registers(0)(244)    <= not(local_tmr_voter(243));                                                                           
                tmr_registers(1)(244)    <= not(local_tmr_voter(243));                                                                           
                tmr_registers(2)(244)    <= not(local_tmr_voter(243));                                                                           
 
                tmr_registers(0)(245)    <= not(local_tmr_voter(244));                                                                           
                tmr_registers(1)(245)    <= not(local_tmr_voter(244));                                                                           
                tmr_registers(2)(245)    <= not(local_tmr_voter(244));                                                                           
 
                tmr_registers(0)(246)    <= not(local_tmr_voter(245));                                                                           
                tmr_registers(1)(246)    <= not(local_tmr_voter(245));                                                                           
                tmr_registers(2)(246)    <= not(local_tmr_voter(245));                                                                           
 
                tmr_registers(0)(247)    <= not(local_tmr_voter(246));                                                                           
                tmr_registers(1)(247)    <= not(local_tmr_voter(246));                                                                           
                tmr_registers(2)(247)    <= not(local_tmr_voter(246));                                                                           
 
                tmr_registers(0)(248)    <= not(local_tmr_voter(247));                                                                           
                tmr_registers(1)(248)    <= not(local_tmr_voter(247));                                                                           
                tmr_registers(2)(248)    <= not(local_tmr_voter(247));                                                                           
 
                tmr_registers(0)(249)    <= not(local_tmr_voter(248));                                                                           
                tmr_registers(1)(249)    <= not(local_tmr_voter(248));                                                                           
                tmr_registers(2)(249)    <= not(local_tmr_voter(248));                                                                           
 
                tmr_registers(0)(250)    <= not(local_tmr_voter(249));                                                                           
                tmr_registers(1)(250)    <= not(local_tmr_voter(249));                                                                           
                tmr_registers(2)(250)    <= not(local_tmr_voter(249));                                                                           
 
                tmr_registers(0)(251)    <= not(local_tmr_voter(250));                                                                           
                tmr_registers(1)(251)    <= not(local_tmr_voter(250));                                                                           
                tmr_registers(2)(251)    <= not(local_tmr_voter(250));                                                                           
 
                tmr_registers(0)(252)    <= not(local_tmr_voter(251));                                                                           
                tmr_registers(1)(252)    <= not(local_tmr_voter(251));                                                                           
                tmr_registers(2)(252)    <= not(local_tmr_voter(251));                                                                           
 
                tmr_registers(0)(253)    <= not(local_tmr_voter(252));                                                                           
                tmr_registers(1)(253)    <= not(local_tmr_voter(252));                                                                           
                tmr_registers(2)(253)    <= not(local_tmr_voter(252));                                                                           
 
                tmr_registers(0)(254)    <= not(local_tmr_voter(253));                                                                           
                tmr_registers(1)(254)    <= not(local_tmr_voter(253));                                                                           
                tmr_registers(2)(254)    <= not(local_tmr_voter(253));                                                                           
 
                tmr_registers(0)(255)    <= not(local_tmr_voter(254));                                                                           
                tmr_registers(1)(255)    <= not(local_tmr_voter(254));                                                                           
                tmr_registers(2)(255)    <= not(local_tmr_voter(254));                                                                           
 
                tmr_registers(0)(256)    <= not(local_tmr_voter(255));                                                                           
                tmr_registers(1)(256)    <= not(local_tmr_voter(255));                                                                           
                tmr_registers(2)(256)    <= not(local_tmr_voter(255));                                                                           
 
                tmr_registers(0)(257)    <= not(local_tmr_voter(256));                                                                           
                tmr_registers(1)(257)    <= not(local_tmr_voter(256));                                                                           
                tmr_registers(2)(257)    <= not(local_tmr_voter(256));                                                                           
 
                tmr_registers(0)(258)    <= not(local_tmr_voter(257));                                                                           
                tmr_registers(1)(258)    <= not(local_tmr_voter(257));                                                                           
                tmr_registers(2)(258)    <= not(local_tmr_voter(257));                                                                           
 
                tmr_registers(0)(259)    <= not(local_tmr_voter(258));                                                                           
                tmr_registers(1)(259)    <= not(local_tmr_voter(258));                                                                           
                tmr_registers(2)(259)    <= not(local_tmr_voter(258));                                                                           
 
                tmr_registers(0)(260)    <= not(local_tmr_voter(259));                                                                           
                tmr_registers(1)(260)    <= not(local_tmr_voter(259));                                                                           
                tmr_registers(2)(260)    <= not(local_tmr_voter(259));                                                                           
 
                tmr_registers(0)(261)    <= not(local_tmr_voter(260));                                                                           
                tmr_registers(1)(261)    <= not(local_tmr_voter(260));                                                                           
                tmr_registers(2)(261)    <= not(local_tmr_voter(260));                                                                           
 
                tmr_registers(0)(262)    <= not(local_tmr_voter(261));                                                                           
                tmr_registers(1)(262)    <= not(local_tmr_voter(261));                                                                           
                tmr_registers(2)(262)    <= not(local_tmr_voter(261));                                                                           
 
                tmr_registers(0)(263)    <= not(local_tmr_voter(262));                                                                           
                tmr_registers(1)(263)    <= not(local_tmr_voter(262));                                                                           
                tmr_registers(2)(263)    <= not(local_tmr_voter(262));                                                                           
 
                tmr_registers(0)(264)    <= not(local_tmr_voter(263));                                                                           
                tmr_registers(1)(264)    <= not(local_tmr_voter(263));                                                                           
                tmr_registers(2)(264)    <= not(local_tmr_voter(263));                                                                           
 
                tmr_registers(0)(265)    <= not(local_tmr_voter(264));                                                                           
                tmr_registers(1)(265)    <= not(local_tmr_voter(264));                                                                           
                tmr_registers(2)(265)    <= not(local_tmr_voter(264));                                                                           
 
                tmr_registers(0)(266)    <= not(local_tmr_voter(265));                                                                           
                tmr_registers(1)(266)    <= not(local_tmr_voter(265));                                                                           
                tmr_registers(2)(266)    <= not(local_tmr_voter(265));                                                                           
 
                tmr_registers(0)(267)    <= not(local_tmr_voter(266));                                                                           
                tmr_registers(1)(267)    <= not(local_tmr_voter(266));                                                                           
                tmr_registers(2)(267)    <= not(local_tmr_voter(266));                                                                           
 
                tmr_registers(0)(268)    <= not(local_tmr_voter(267));                                                                           
                tmr_registers(1)(268)    <= not(local_tmr_voter(267));                                                                           
                tmr_registers(2)(268)    <= not(local_tmr_voter(267));                                                                           
 
                tmr_registers(0)(269)    <= not(local_tmr_voter(268));                                                                           
                tmr_registers(1)(269)    <= not(local_tmr_voter(268));                                                                           
                tmr_registers(2)(269)    <= not(local_tmr_voter(268));                                                                           
 
                tmr_registers(0)(270)    <= not(local_tmr_voter(269));                                                                           
                tmr_registers(1)(270)    <= not(local_tmr_voter(269));                                                                           
                tmr_registers(2)(270)    <= not(local_tmr_voter(269));                                                                           
 
                tmr_registers(0)(271)    <= not(local_tmr_voter(270));                                                                           
                tmr_registers(1)(271)    <= not(local_tmr_voter(270));                                                                           
                tmr_registers(2)(271)    <= not(local_tmr_voter(270));                                                                           
 
                tmr_registers(0)(272)    <= not(local_tmr_voter(271));                                                                           
                tmr_registers(1)(272)    <= not(local_tmr_voter(271));                                                                           
                tmr_registers(2)(272)    <= not(local_tmr_voter(271));                                                                           
 
                tmr_registers(0)(273)    <= not(local_tmr_voter(272));                                                                           
                tmr_registers(1)(273)    <= not(local_tmr_voter(272));                                                                           
                tmr_registers(2)(273)    <= not(local_tmr_voter(272));                                                                           
 
                tmr_registers(0)(274)    <= not(local_tmr_voter(273));                                                                           
                tmr_registers(1)(274)    <= not(local_tmr_voter(273));                                                                           
                tmr_registers(2)(274)    <= not(local_tmr_voter(273));                                                                           
 
                tmr_registers(0)(275)    <= not(local_tmr_voter(274));                                                                           
                tmr_registers(1)(275)    <= not(local_tmr_voter(274));                                                                           
                tmr_registers(2)(275)    <= not(local_tmr_voter(274));                                                                           
 
                tmr_registers(0)(276)    <= not(local_tmr_voter(275));                                                                           
                tmr_registers(1)(276)    <= not(local_tmr_voter(275));                                                                           
                tmr_registers(2)(276)    <= not(local_tmr_voter(275));                                                                           
 
                tmr_registers(0)(277)    <= not(local_tmr_voter(276));                                                                           
                tmr_registers(1)(277)    <= not(local_tmr_voter(276));                                                                           
                tmr_registers(2)(277)    <= not(local_tmr_voter(276));                                                                           
 
                tmr_registers(0)(278)    <= not(local_tmr_voter(277));                                                                           
                tmr_registers(1)(278)    <= not(local_tmr_voter(277));                                                                           
                tmr_registers(2)(278)    <= not(local_tmr_voter(277));                                                                           
 
                tmr_registers(0)(279)    <= not(local_tmr_voter(278));                                                                           
                tmr_registers(1)(279)    <= not(local_tmr_voter(278));                                                                           
                tmr_registers(2)(279)    <= not(local_tmr_voter(278));                                                                           
 
                tmr_registers(0)(280)    <= not(local_tmr_voter(279));                                                                           
                tmr_registers(1)(280)    <= not(local_tmr_voter(279));                                                                           
                tmr_registers(2)(280)    <= not(local_tmr_voter(279));                                                                           
 
                tmr_registers(0)(281)    <= not(local_tmr_voter(280));                                                                           
                tmr_registers(1)(281)    <= not(local_tmr_voter(280));                                                                           
                tmr_registers(2)(281)    <= not(local_tmr_voter(280));                                                                           
 
                tmr_registers(0)(282)    <= not(local_tmr_voter(281));                                                                           
                tmr_registers(1)(282)    <= not(local_tmr_voter(281));                                                                           
                tmr_registers(2)(282)    <= not(local_tmr_voter(281));                                                                           
 
                tmr_registers(0)(283)    <= not(local_tmr_voter(282));                                                                           
                tmr_registers(1)(283)    <= not(local_tmr_voter(282));                                                                           
                tmr_registers(2)(283)    <= not(local_tmr_voter(282));                                                                           
 
                tmr_registers(0)(284)    <= not(local_tmr_voter(283));                                                                           
                tmr_registers(1)(284)    <= not(local_tmr_voter(283));                                                                           
                tmr_registers(2)(284)    <= not(local_tmr_voter(283));                                                                           
 
                tmr_registers(0)(285)    <= not(local_tmr_voter(284));                                                                           
                tmr_registers(1)(285)    <= not(local_tmr_voter(284));                                                                           
                tmr_registers(2)(285)    <= not(local_tmr_voter(284));                                                                           
 
                tmr_registers(0)(286)    <= not(local_tmr_voter(285));                                                                           
                tmr_registers(1)(286)    <= not(local_tmr_voter(285));                                                                           
                tmr_registers(2)(286)    <= not(local_tmr_voter(285));                                                                           
 
                tmr_registers(0)(287)    <= not(local_tmr_voter(286));                                                                           
                tmr_registers(1)(287)    <= not(local_tmr_voter(286));                                                                           
                tmr_registers(2)(287)    <= not(local_tmr_voter(286));                                                                           
 
                tmr_registers(0)(288)    <= not(local_tmr_voter(287));                                                                           
                tmr_registers(1)(288)    <= not(local_tmr_voter(287));                                                                           
                tmr_registers(2)(288)    <= not(local_tmr_voter(287));                                                                           
 
                tmr_registers(0)(289)    <= not(local_tmr_voter(288));                                                                           
                tmr_registers(1)(289)    <= not(local_tmr_voter(288));                                                                           
                tmr_registers(2)(289)    <= not(local_tmr_voter(288));                                                                           
 
                tmr_registers(0)(290)    <= not(local_tmr_voter(289));                                                                           
                tmr_registers(1)(290)    <= not(local_tmr_voter(289));                                                                           
                tmr_registers(2)(290)    <= not(local_tmr_voter(289));                                                                           
 
                tmr_registers(0)(291)    <= not(local_tmr_voter(290));                                                                           
                tmr_registers(1)(291)    <= not(local_tmr_voter(290));                                                                           
                tmr_registers(2)(291)    <= not(local_tmr_voter(290));                                                                           
 
                tmr_registers(0)(292)    <= not(local_tmr_voter(291));                                                                           
                tmr_registers(1)(292)    <= not(local_tmr_voter(291));                                                                           
                tmr_registers(2)(292)    <= not(local_tmr_voter(291));                                                                           
 
                tmr_registers(0)(293)    <= not(local_tmr_voter(292));                                                                           
                tmr_registers(1)(293)    <= not(local_tmr_voter(292));                                                                           
                tmr_registers(2)(293)    <= not(local_tmr_voter(292));                                                                           
 
                tmr_registers(0)(294)    <= not(local_tmr_voter(293));                                                                           
                tmr_registers(1)(294)    <= not(local_tmr_voter(293));                                                                           
                tmr_registers(2)(294)    <= not(local_tmr_voter(293));                                                                           
 
                tmr_registers(0)(295)    <= not(local_tmr_voter(294));                                                                           
                tmr_registers(1)(295)    <= not(local_tmr_voter(294));                                                                           
                tmr_registers(2)(295)    <= not(local_tmr_voter(294));                                                                           
 
                tmr_registers(0)(296)    <= not(local_tmr_voter(295));                                                                           
                tmr_registers(1)(296)    <= not(local_tmr_voter(295));                                                                           
                tmr_registers(2)(296)    <= not(local_tmr_voter(295));                                                                           
 
                tmr_registers(0)(297)    <= not(local_tmr_voter(296));                                                                           
                tmr_registers(1)(297)    <= not(local_tmr_voter(296));                                                                           
                tmr_registers(2)(297)    <= not(local_tmr_voter(296));                                                                           
 
                tmr_registers(0)(298)    <= not(local_tmr_voter(297));                                                                           
                tmr_registers(1)(298)    <= not(local_tmr_voter(297));                                                                           
                tmr_registers(2)(298)    <= not(local_tmr_voter(297));                                                                           
 
                tmr_registers(0)(299)    <= not(local_tmr_voter(298));                                                                           
                tmr_registers(1)(299)    <= not(local_tmr_voter(298));                                                                           
                tmr_registers(2)(299)    <= not(local_tmr_voter(298));                                                                           
 
                tmr_registers(0)(300)    <= not(local_tmr_voter(299));                                                                           
                tmr_registers(1)(300)    <= not(local_tmr_voter(299));                                                                           
                tmr_registers(2)(300)    <= not(local_tmr_voter(299));                                                                           
 
                tmr_registers(0)(301)    <= not(local_tmr_voter(300));                                                                           
                tmr_registers(1)(301)    <= not(local_tmr_voter(300));                                                                           
                tmr_registers(2)(301)    <= not(local_tmr_voter(300));                                                                           
 
                tmr_registers(0)(302)    <= not(local_tmr_voter(301));                                                                           
                tmr_registers(1)(302)    <= not(local_tmr_voter(301));                                                                           
                tmr_registers(2)(302)    <= not(local_tmr_voter(301));                                                                           
 
                tmr_registers(0)(303)    <= not(local_tmr_voter(302));                                                                           
                tmr_registers(1)(303)    <= not(local_tmr_voter(302));                                                                           
                tmr_registers(2)(303)    <= not(local_tmr_voter(302));                                                                           
 
                tmr_registers(0)(304)    <= not(local_tmr_voter(303));                                                                           
                tmr_registers(1)(304)    <= not(local_tmr_voter(303));                                                                           
                tmr_registers(2)(304)    <= not(local_tmr_voter(303));                                                                           
 
                tmr_registers(0)(305)    <= not(local_tmr_voter(304));                                                                           
                tmr_registers(1)(305)    <= not(local_tmr_voter(304));                                                                           
                tmr_registers(2)(305)    <= not(local_tmr_voter(304));                                                                           
 
                tmr_registers(0)(306)    <= not(local_tmr_voter(305));                                                                           
                tmr_registers(1)(306)    <= not(local_tmr_voter(305));                                                                           
                tmr_registers(2)(306)    <= not(local_tmr_voter(305));                                                                           
 
                tmr_registers(0)(307)    <= not(local_tmr_voter(306));                                                                           
                tmr_registers(1)(307)    <= not(local_tmr_voter(306));                                                                           
                tmr_registers(2)(307)    <= not(local_tmr_voter(306));                                                                           
 
                tmr_registers(0)(308)    <= not(local_tmr_voter(307));                                                                           
                tmr_registers(1)(308)    <= not(local_tmr_voter(307));                                                                           
                tmr_registers(2)(308)    <= not(local_tmr_voter(307));                                                                           
 
                tmr_registers(0)(309)    <= not(local_tmr_voter(308));                                                                           
                tmr_registers(1)(309)    <= not(local_tmr_voter(308));                                                                           
                tmr_registers(2)(309)    <= not(local_tmr_voter(308));                                                                           
 
                tmr_registers(0)(310)    <= not(local_tmr_voter(309));                                                                           
                tmr_registers(1)(310)    <= not(local_tmr_voter(309));                                                                           
                tmr_registers(2)(310)    <= not(local_tmr_voter(309));                                                                           
 
                tmr_registers(0)(311)    <= not(local_tmr_voter(310));                                                                           
                tmr_registers(1)(311)    <= not(local_tmr_voter(310));                                                                           
                tmr_registers(2)(311)    <= not(local_tmr_voter(310));                                                                           
 
                tmr_registers(0)(312)    <= not(local_tmr_voter(311));                                                                           
                tmr_registers(1)(312)    <= not(local_tmr_voter(311));                                                                           
                tmr_registers(2)(312)    <= not(local_tmr_voter(311));                                                                           
 
                tmr_registers(0)(313)    <= not(local_tmr_voter(312));                                                                           
                tmr_registers(1)(313)    <= not(local_tmr_voter(312));                                                                           
                tmr_registers(2)(313)    <= not(local_tmr_voter(312));                                                                           
 
                tmr_registers(0)(314)    <= not(local_tmr_voter(313));                                                                           
                tmr_registers(1)(314)    <= not(local_tmr_voter(313));                                                                           
                tmr_registers(2)(314)    <= not(local_tmr_voter(313));                                                                           
 
                tmr_registers(0)(315)    <= not(local_tmr_voter(314));                                                                           
                tmr_registers(1)(315)    <= not(local_tmr_voter(314));                                                                           
                tmr_registers(2)(315)    <= not(local_tmr_voter(314));                                                                           
 
                tmr_registers(0)(316)    <= not(local_tmr_voter(315));                                                                           
                tmr_registers(1)(316)    <= not(local_tmr_voter(315));                                                                           
                tmr_registers(2)(316)    <= not(local_tmr_voter(315));                                                                           
 
                tmr_registers(0)(317)    <= not(local_tmr_voter(316));                                                                           
                tmr_registers(1)(317)    <= not(local_tmr_voter(316));                                                                           
                tmr_registers(2)(317)    <= not(local_tmr_voter(316));                                                                           
 
                tmr_registers(0)(318)    <= not(local_tmr_voter(317));                                                                           
                tmr_registers(1)(318)    <= not(local_tmr_voter(317));                                                                           
                tmr_registers(2)(318)    <= not(local_tmr_voter(317));                                                                           
 
                tmr_registers(0)(319)    <= not(local_tmr_voter(318));                                                                           
                tmr_registers(1)(319)    <= not(local_tmr_voter(318));                                                                           
                tmr_registers(2)(319)    <= not(local_tmr_voter(318));                                                                           
 
                tmr_registers(0)(320)    <= not(local_tmr_voter(319));                                                                           
                tmr_registers(1)(320)    <= not(local_tmr_voter(319));                                                                           
                tmr_registers(2)(320)    <= not(local_tmr_voter(319));                                                                           
 
                tmr_registers(0)(321)    <= not(local_tmr_voter(320));                                                                           
                tmr_registers(1)(321)    <= not(local_tmr_voter(320));                                                                           
                tmr_registers(2)(321)    <= not(local_tmr_voter(320));                                                                           
 
                tmr_registers(0)(322)    <= not(local_tmr_voter(321));                                                                           
                tmr_registers(1)(322)    <= not(local_tmr_voter(321));                                                                           
                tmr_registers(2)(322)    <= not(local_tmr_voter(321));                                                                           
 
                tmr_registers(0)(323)    <= not(local_tmr_voter(322));                                                                           
                tmr_registers(1)(323)    <= not(local_tmr_voter(322));                                                                           
                tmr_registers(2)(323)    <= not(local_tmr_voter(322));                                                                           
 
                tmr_registers(0)(324)    <= not(local_tmr_voter(323));                                                                           
                tmr_registers(1)(324)    <= not(local_tmr_voter(323));                                                                           
                tmr_registers(2)(324)    <= not(local_tmr_voter(323));                                                                           
 
                tmr_registers(0)(325)    <= not(local_tmr_voter(324));                                                                           
                tmr_registers(1)(325)    <= not(local_tmr_voter(324));                                                                           
                tmr_registers(2)(325)    <= not(local_tmr_voter(324));                                                                           
 
                tmr_registers(0)(326)    <= not(local_tmr_voter(325));                                                                           
                tmr_registers(1)(326)    <= not(local_tmr_voter(325));                                                                           
                tmr_registers(2)(326)    <= not(local_tmr_voter(325));                                                                           
 
                tmr_registers(0)(327)    <= not(local_tmr_voter(326));                                                                           
                tmr_registers(1)(327)    <= not(local_tmr_voter(326));                                                                           
                tmr_registers(2)(327)    <= not(local_tmr_voter(326));                                                                           
 
                tmr_registers(0)(328)    <= not(local_tmr_voter(327));                                                                           
                tmr_registers(1)(328)    <= not(local_tmr_voter(327));                                                                           
                tmr_registers(2)(328)    <= not(local_tmr_voter(327));                                                                           
 
                tmr_registers(0)(329)    <= not(local_tmr_voter(328));                                                                           
                tmr_registers(1)(329)    <= not(local_tmr_voter(328));                                                                           
                tmr_registers(2)(329)    <= not(local_tmr_voter(328));                                                                           
 
                tmr_registers(0)(330)    <= not(local_tmr_voter(329));                                                                           
                tmr_registers(1)(330)    <= not(local_tmr_voter(329));                                                                           
                tmr_registers(2)(330)    <= not(local_tmr_voter(329));                                                                           
 
                tmr_registers(0)(331)    <= not(local_tmr_voter(330));                                                                           
                tmr_registers(1)(331)    <= not(local_tmr_voter(330));                                                                           
                tmr_registers(2)(331)    <= not(local_tmr_voter(330));                                                                           
 
                tmr_registers(0)(332)    <= not(local_tmr_voter(331));                                                                           
                tmr_registers(1)(332)    <= not(local_tmr_voter(331));                                                                           
                tmr_registers(2)(332)    <= not(local_tmr_voter(331));                                                                           
 
                tmr_registers(0)(333)    <= not(local_tmr_voter(332));                                                                           
                tmr_registers(1)(333)    <= not(local_tmr_voter(332));                                                                           
                tmr_registers(2)(333)    <= not(local_tmr_voter(332));                                                                           
 
                tmr_registers(0)(334)    <= not(local_tmr_voter(333));                                                                           
                tmr_registers(1)(334)    <= not(local_tmr_voter(333));                                                                           
                tmr_registers(2)(334)    <= not(local_tmr_voter(333));                                                                           
 
                tmr_registers(0)(335)    <= not(local_tmr_voter(334));                                                                           
                tmr_registers(1)(335)    <= not(local_tmr_voter(334));                                                                           
                tmr_registers(2)(335)    <= not(local_tmr_voter(334));                                                                           
 
                tmr_registers(0)(336)    <= not(local_tmr_voter(335));                                                                           
                tmr_registers(1)(336)    <= not(local_tmr_voter(335));                                                                           
                tmr_registers(2)(336)    <= not(local_tmr_voter(335));                                                                           
 
                tmr_registers(0)(337)    <= not(local_tmr_voter(336));                                                                           
                tmr_registers(1)(337)    <= not(local_tmr_voter(336));                                                                           
                tmr_registers(2)(337)    <= not(local_tmr_voter(336));                                                                           
 
                tmr_registers(0)(338)    <= not(local_tmr_voter(337));                                                                           
                tmr_registers(1)(338)    <= not(local_tmr_voter(337));                                                                           
                tmr_registers(2)(338)    <= not(local_tmr_voter(337));                                                                           
 
                tmr_registers(0)(339)    <= not(local_tmr_voter(338));                                                                           
                tmr_registers(1)(339)    <= not(local_tmr_voter(338));                                                                           
                tmr_registers(2)(339)    <= not(local_tmr_voter(338));                                                                           
 
                tmr_registers(0)(340)    <= not(local_tmr_voter(339));                                                                           
                tmr_registers(1)(340)    <= not(local_tmr_voter(339));                                                                           
                tmr_registers(2)(340)    <= not(local_tmr_voter(339));                                                                           
 
                tmr_registers(0)(341)    <= not(local_tmr_voter(340));                                                                           
                tmr_registers(1)(341)    <= not(local_tmr_voter(340));                                                                           
                tmr_registers(2)(341)    <= not(local_tmr_voter(340));                                                                           
 
                tmr_registers(0)(342)    <= not(local_tmr_voter(341));                                                                           
                tmr_registers(1)(342)    <= not(local_tmr_voter(341));                                                                           
                tmr_registers(2)(342)    <= not(local_tmr_voter(341));                                                                           
 
                tmr_registers(0)(343)    <= not(local_tmr_voter(342));                                                                           
                tmr_registers(1)(343)    <= not(local_tmr_voter(342));                                                                           
                tmr_registers(2)(343)    <= not(local_tmr_voter(342));                                                                           
 
                tmr_registers(0)(344)    <= not(local_tmr_voter(343));                                                                           
                tmr_registers(1)(344)    <= not(local_tmr_voter(343));                                                                           
                tmr_registers(2)(344)    <= not(local_tmr_voter(343));                                                                           
 
                tmr_registers(0)(345)    <= not(local_tmr_voter(344));                                                                           
                tmr_registers(1)(345)    <= not(local_tmr_voter(344));                                                                           
                tmr_registers(2)(345)    <= not(local_tmr_voter(344));                                                                           
 
                tmr_registers(0)(346)    <= not(local_tmr_voter(345));                                                                           
                tmr_registers(1)(346)    <= not(local_tmr_voter(345));                                                                           
                tmr_registers(2)(346)    <= not(local_tmr_voter(345));                                                                           
 
                tmr_registers(0)(347)    <= not(local_tmr_voter(346));                                                                           
                tmr_registers(1)(347)    <= not(local_tmr_voter(346));                                                                           
                tmr_registers(2)(347)    <= not(local_tmr_voter(346));                                                                           
 
                tmr_registers(0)(348)    <= not(local_tmr_voter(347));                                                                           
                tmr_registers(1)(348)    <= not(local_tmr_voter(347));                                                                           
                tmr_registers(2)(348)    <= not(local_tmr_voter(347));                                                                           
 
                tmr_registers(0)(349)    <= not(local_tmr_voter(348));                                                                           
                tmr_registers(1)(349)    <= not(local_tmr_voter(348));                                                                           
                tmr_registers(2)(349)    <= not(local_tmr_voter(348));                                                                           
 
                tmr_registers(0)(350)    <= not(local_tmr_voter(349));                                                                           
                tmr_registers(1)(350)    <= not(local_tmr_voter(349));                                                                           
                tmr_registers(2)(350)    <= not(local_tmr_voter(349));                                                                           
 
                tmr_registers(0)(351)    <= not(local_tmr_voter(350));                                                                           
                tmr_registers(1)(351)    <= not(local_tmr_voter(350));                                                                           
                tmr_registers(2)(351)    <= not(local_tmr_voter(350));                                                                           
 
                tmr_registers(0)(352)    <= not(local_tmr_voter(351));                                                                           
                tmr_registers(1)(352)    <= not(local_tmr_voter(351));                                                                           
                tmr_registers(2)(352)    <= not(local_tmr_voter(351));                                                                           
 
                tmr_registers(0)(353)    <= not(local_tmr_voter(352));                                                                           
                tmr_registers(1)(353)    <= not(local_tmr_voter(352));                                                                           
                tmr_registers(2)(353)    <= not(local_tmr_voter(352));                                                                           
 
                tmr_registers(0)(354)    <= not(local_tmr_voter(353));                                                                           
                tmr_registers(1)(354)    <= not(local_tmr_voter(353));                                                                           
                tmr_registers(2)(354)    <= not(local_tmr_voter(353));                                                                           
 
                tmr_registers(0)(355)    <= not(local_tmr_voter(354));                                                                           
                tmr_registers(1)(355)    <= not(local_tmr_voter(354));                                                                           
                tmr_registers(2)(355)    <= not(local_tmr_voter(354));                                                                           
 
                tmr_registers(0)(356)    <= not(local_tmr_voter(355));                                                                           
                tmr_registers(1)(356)    <= not(local_tmr_voter(355));                                                                           
                tmr_registers(2)(356)    <= not(local_tmr_voter(355));                                                                           
 
                tmr_registers(0)(357)    <= not(local_tmr_voter(356));                                                                           
                tmr_registers(1)(357)    <= not(local_tmr_voter(356));                                                                           
                tmr_registers(2)(357)    <= not(local_tmr_voter(356));                                                                           
 
                tmr_registers(0)(358)    <= not(local_tmr_voter(357));                                                                           
                tmr_registers(1)(358)    <= not(local_tmr_voter(357));                                                                           
                tmr_registers(2)(358)    <= not(local_tmr_voter(357));                                                                           
 
                tmr_registers(0)(359)    <= not(local_tmr_voter(358));                                                                           
                tmr_registers(1)(359)    <= not(local_tmr_voter(358));                                                                           
                tmr_registers(2)(359)    <= not(local_tmr_voter(358));                                                                           
 
                tmr_registers(0)(360)    <= not(local_tmr_voter(359));                                                                           
                tmr_registers(1)(360)    <= not(local_tmr_voter(359));                                                                           
                tmr_registers(2)(360)    <= not(local_tmr_voter(359));                                                                           
 
                tmr_registers(0)(361)    <= not(local_tmr_voter(360));                                                                           
                tmr_registers(1)(361)    <= not(local_tmr_voter(360));                                                                           
                tmr_registers(2)(361)    <= not(local_tmr_voter(360));                                                                           
 
                tmr_registers(0)(362)    <= not(local_tmr_voter(361));                                                                           
                tmr_registers(1)(362)    <= not(local_tmr_voter(361));                                                                           
                tmr_registers(2)(362)    <= not(local_tmr_voter(361));                                                                           
 
                tmr_registers(0)(363)    <= not(local_tmr_voter(362));                                                                           
                tmr_registers(1)(363)    <= not(local_tmr_voter(362));                                                                           
                tmr_registers(2)(363)    <= not(local_tmr_voter(362));                                                                           
 
                tmr_registers(0)(364)    <= not(local_tmr_voter(363));                                                                           
                tmr_registers(1)(364)    <= not(local_tmr_voter(363));                                                                           
                tmr_registers(2)(364)    <= not(local_tmr_voter(363));                                                                           
 
                tmr_registers(0)(365)    <= not(local_tmr_voter(364));                                                                           
                tmr_registers(1)(365)    <= not(local_tmr_voter(364));                                                                           
                tmr_registers(2)(365)    <= not(local_tmr_voter(364));                                                                           
 
                tmr_registers(0)(366)    <= not(local_tmr_voter(365));                                                                           
                tmr_registers(1)(366)    <= not(local_tmr_voter(365));                                                                           
                tmr_registers(2)(366)    <= not(local_tmr_voter(365));                                                                           
 
                tmr_registers(0)(367)    <= not(local_tmr_voter(366));                                                                           
                tmr_registers(1)(367)    <= not(local_tmr_voter(366));                                                                           
                tmr_registers(2)(367)    <= not(local_tmr_voter(366));                                                                           
 
                tmr_registers(0)(368)    <= not(local_tmr_voter(367));                                                                           
                tmr_registers(1)(368)    <= not(local_tmr_voter(367));                                                                           
                tmr_registers(2)(368)    <= not(local_tmr_voter(367));                                                                           
 
                tmr_registers(0)(369)    <= not(local_tmr_voter(368));                                                                           
                tmr_registers(1)(369)    <= not(local_tmr_voter(368));                                                                           
                tmr_registers(2)(369)    <= not(local_tmr_voter(368));                                                                           
 
                tmr_registers(0)(370)    <= not(local_tmr_voter(369));                                                                           
                tmr_registers(1)(370)    <= not(local_tmr_voter(369));                                                                           
                tmr_registers(2)(370)    <= not(local_tmr_voter(369));                                                                           
 
                tmr_registers(0)(371)    <= not(local_tmr_voter(370));                                                                           
                tmr_registers(1)(371)    <= not(local_tmr_voter(370));                                                                           
                tmr_registers(2)(371)    <= not(local_tmr_voter(370));                                                                           
 
                tmr_registers(0)(372)    <= not(local_tmr_voter(371));                                                                           
                tmr_registers(1)(372)    <= not(local_tmr_voter(371));                                                                           
                tmr_registers(2)(372)    <= not(local_tmr_voter(371));                                                                           
 
                tmr_registers(0)(373)    <= not(local_tmr_voter(372));                                                                           
                tmr_registers(1)(373)    <= not(local_tmr_voter(372));                                                                           
                tmr_registers(2)(373)    <= not(local_tmr_voter(372));                                                                           
 
                tmr_registers(0)(374)    <= not(local_tmr_voter(373));                                                                           
                tmr_registers(1)(374)    <= not(local_tmr_voter(373));                                                                           
                tmr_registers(2)(374)    <= not(local_tmr_voter(373));                                                                           
 
                tmr_registers(0)(375)    <= not(local_tmr_voter(374));                                                                           
                tmr_registers(1)(375)    <= not(local_tmr_voter(374));                                                                           
                tmr_registers(2)(375)    <= not(local_tmr_voter(374));                                                                           
 
                tmr_registers(0)(376)    <= not(local_tmr_voter(375));                                                                           
                tmr_registers(1)(376)    <= not(local_tmr_voter(375));                                                                           
                tmr_registers(2)(376)    <= not(local_tmr_voter(375));                                                                           
 
                tmr_registers(0)(377)    <= not(local_tmr_voter(376));                                                                           
                tmr_registers(1)(377)    <= not(local_tmr_voter(376));                                                                           
                tmr_registers(2)(377)    <= not(local_tmr_voter(376));                                                                           
 
                tmr_registers(0)(378)    <= not(local_tmr_voter(377));                                                                           
                tmr_registers(1)(378)    <= not(local_tmr_voter(377));                                                                           
                tmr_registers(2)(378)    <= not(local_tmr_voter(377));                                                                           
 
                tmr_registers(0)(379)    <= not(local_tmr_voter(378));                                                                           
                tmr_registers(1)(379)    <= not(local_tmr_voter(378));                                                                           
                tmr_registers(2)(379)    <= not(local_tmr_voter(378));                                                                           
 
                tmr_registers(0)(380)    <= not(local_tmr_voter(379));                                                                           
                tmr_registers(1)(380)    <= not(local_tmr_voter(379));                                                                           
                tmr_registers(2)(380)    <= not(local_tmr_voter(379));                                                                           
 
                tmr_registers(0)(381)    <= not(local_tmr_voter(380));                                                                           
                tmr_registers(1)(381)    <= not(local_tmr_voter(380));                                                                           
                tmr_registers(2)(381)    <= not(local_tmr_voter(380));                                                                           
 
                tmr_registers(0)(382)    <= not(local_tmr_voter(381));                                                                           
                tmr_registers(1)(382)    <= not(local_tmr_voter(381));                                                                           
                tmr_registers(2)(382)    <= not(local_tmr_voter(381));                                                                           
 
                tmr_registers(0)(383)    <= not(local_tmr_voter(382));                                                                           
                tmr_registers(1)(383)    <= not(local_tmr_voter(382));                                                                           
                tmr_registers(2)(383)    <= not(local_tmr_voter(382));                                                                           
 
                tmr_registers(0)(384)    <= not(local_tmr_voter(383));                                                                           
                tmr_registers(1)(384)    <= not(local_tmr_voter(383));                                                                           
                tmr_registers(2)(384)    <= not(local_tmr_voter(383));                                                                           
 
                tmr_registers(0)(385)    <= not(local_tmr_voter(384));                                                                           
                tmr_registers(1)(385)    <= not(local_tmr_voter(384));                                                                           
                tmr_registers(2)(385)    <= not(local_tmr_voter(384));                                                                           
 
                tmr_registers(0)(386)    <= not(local_tmr_voter(385));                                                                           
                tmr_registers(1)(386)    <= not(local_tmr_voter(385));                                                                           
                tmr_registers(2)(386)    <= not(local_tmr_voter(385));                                                                           
 
                tmr_registers(0)(387)    <= not(local_tmr_voter(386));                                                                           
                tmr_registers(1)(387)    <= not(local_tmr_voter(386));                                                                           
                tmr_registers(2)(387)    <= not(local_tmr_voter(386));                                                                           
 
                tmr_registers(0)(388)    <= not(local_tmr_voter(387));                                                                           
                tmr_registers(1)(388)    <= not(local_tmr_voter(387));                                                                           
                tmr_registers(2)(388)    <= not(local_tmr_voter(387));                                                                           
 
                tmr_registers(0)(389)    <= not(local_tmr_voter(388));                                                                           
                tmr_registers(1)(389)    <= not(local_tmr_voter(388));                                                                           
                tmr_registers(2)(389)    <= not(local_tmr_voter(388));                                                                           
 
                tmr_registers(0)(390)    <= not(local_tmr_voter(389));                                                                           
                tmr_registers(1)(390)    <= not(local_tmr_voter(389));                                                                           
                tmr_registers(2)(390)    <= not(local_tmr_voter(389));                                                                           
 
                tmr_registers(0)(391)    <= not(local_tmr_voter(390));                                                                           
                tmr_registers(1)(391)    <= not(local_tmr_voter(390));                                                                           
                tmr_registers(2)(391)    <= not(local_tmr_voter(390));                                                                           
 
                tmr_registers(0)(392)    <= not(local_tmr_voter(391));                                                                           
                tmr_registers(1)(392)    <= not(local_tmr_voter(391));                                                                           
                tmr_registers(2)(392)    <= not(local_tmr_voter(391));                                                                           
 
                tmr_registers(0)(393)    <= not(local_tmr_voter(392));                                                                           
                tmr_registers(1)(393)    <= not(local_tmr_voter(392));                                                                           
                tmr_registers(2)(393)    <= not(local_tmr_voter(392));                                                                           
 
                tmr_registers(0)(394)    <= not(local_tmr_voter(393));                                                                           
                tmr_registers(1)(394)    <= not(local_tmr_voter(393));                                                                           
                tmr_registers(2)(394)    <= not(local_tmr_voter(393));                                                                           
 
                tmr_registers(0)(395)    <= not(local_tmr_voter(394));                                                                           
                tmr_registers(1)(395)    <= not(local_tmr_voter(394));                                                                           
                tmr_registers(2)(395)    <= not(local_tmr_voter(394));                                                                           
 
                tmr_registers(0)(396)    <= not(local_tmr_voter(395));                                                                           
                tmr_registers(1)(396)    <= not(local_tmr_voter(395));                                                                           
                tmr_registers(2)(396)    <= not(local_tmr_voter(395));                                                                           
 
                tmr_registers(0)(397)    <= not(local_tmr_voter(396));                                                                           
                tmr_registers(1)(397)    <= not(local_tmr_voter(396));                                                                           
                tmr_registers(2)(397)    <= not(local_tmr_voter(396));                                                                           
 
                tmr_registers(0)(398)    <= not(local_tmr_voter(397));                                                                           
                tmr_registers(1)(398)    <= not(local_tmr_voter(397));                                                                           
                tmr_registers(2)(398)    <= not(local_tmr_voter(397));                                                                           
 
                tmr_registers(0)(399)    <= not(local_tmr_voter(398));                                                                           
                tmr_registers(1)(399)    <= not(local_tmr_voter(398));                                                                           
                tmr_registers(2)(399)    <= not(local_tmr_voter(398));                                                                           
 
                tmr_registers(0)(400)    <= not(local_tmr_voter(399));                                                                           
                tmr_registers(1)(400)    <= not(local_tmr_voter(399));                                                                           
                tmr_registers(2)(400)    <= not(local_tmr_voter(399));                                                                           
 
                tmr_registers(0)(401)    <= not(local_tmr_voter(400));                                                                           
                tmr_registers(1)(401)    <= not(local_tmr_voter(400));                                                                           
                tmr_registers(2)(401)    <= not(local_tmr_voter(400));                                                                           
 
                tmr_registers(0)(402)    <= not(local_tmr_voter(401));                                                                           
                tmr_registers(1)(402)    <= not(local_tmr_voter(401));                                                                           
                tmr_registers(2)(402)    <= not(local_tmr_voter(401));                                                                           
 
                tmr_registers(0)(403)    <= not(local_tmr_voter(402));                                                                           
                tmr_registers(1)(403)    <= not(local_tmr_voter(402));                                                                           
                tmr_registers(2)(403)    <= not(local_tmr_voter(402));                                                                           
 
                tmr_registers(0)(404)    <= not(local_tmr_voter(403));                                                                           
                tmr_registers(1)(404)    <= not(local_tmr_voter(403));                                                                           
                tmr_registers(2)(404)    <= not(local_tmr_voter(403));                                                                           
 
                tmr_registers(0)(405)    <= not(local_tmr_voter(404));                                                                           
                tmr_registers(1)(405)    <= not(local_tmr_voter(404));                                                                           
                tmr_registers(2)(405)    <= not(local_tmr_voter(404));                                                                           
 
                tmr_registers(0)(406)    <= not(local_tmr_voter(405));                                                                           
                tmr_registers(1)(406)    <= not(local_tmr_voter(405));                                                                           
                tmr_registers(2)(406)    <= not(local_tmr_voter(405));                                                                           
 
                tmr_registers(0)(407)    <= not(local_tmr_voter(406));                                                                           
                tmr_registers(1)(407)    <= not(local_tmr_voter(406));                                                                           
                tmr_registers(2)(407)    <= not(local_tmr_voter(406));                                                                           
 
                tmr_registers(0)(408)    <= not(local_tmr_voter(407));                                                                           
                tmr_registers(1)(408)    <= not(local_tmr_voter(407));                                                                           
                tmr_registers(2)(408)    <= not(local_tmr_voter(407));                                                                           
 
                tmr_registers(0)(409)    <= not(local_tmr_voter(408));                                                                           
                tmr_registers(1)(409)    <= not(local_tmr_voter(408));                                                                           
                tmr_registers(2)(409)    <= not(local_tmr_voter(408));                                                                           
 
                tmr_registers(0)(410)    <= not(local_tmr_voter(409));                                                                           
                tmr_registers(1)(410)    <= not(local_tmr_voter(409));                                                                           
                tmr_registers(2)(410)    <= not(local_tmr_voter(409));                                                                           
 
                tmr_registers(0)(411)    <= not(local_tmr_voter(410));                                                                           
                tmr_registers(1)(411)    <= not(local_tmr_voter(410));                                                                           
                tmr_registers(2)(411)    <= not(local_tmr_voter(410));                                                                           
 
                tmr_registers(0)(412)    <= not(local_tmr_voter(411));                                                                           
                tmr_registers(1)(412)    <= not(local_tmr_voter(411));                                                                           
                tmr_registers(2)(412)    <= not(local_tmr_voter(411));                                                                           
 
                tmr_registers(0)(413)    <= not(local_tmr_voter(412));                                                                           
                tmr_registers(1)(413)    <= not(local_tmr_voter(412));                                                                           
                tmr_registers(2)(413)    <= not(local_tmr_voter(412));                                                                           
 
                tmr_registers(0)(414)    <= not(local_tmr_voter(413));                                                                           
                tmr_registers(1)(414)    <= not(local_tmr_voter(413));                                                                           
                tmr_registers(2)(414)    <= not(local_tmr_voter(413));                                                                           
 
                tmr_registers(0)(415)    <= not(local_tmr_voter(414));                                                                           
                tmr_registers(1)(415)    <= not(local_tmr_voter(414));                                                                           
                tmr_registers(2)(415)    <= not(local_tmr_voter(414));                                                                           
 
                tmr_registers(0)(416)    <= not(local_tmr_voter(415));                                                                           
                tmr_registers(1)(416)    <= not(local_tmr_voter(415));                                                                           
                tmr_registers(2)(416)    <= not(local_tmr_voter(415));                                                                           
 
                tmr_registers(0)(417)    <= not(local_tmr_voter(416));                                                                           
                tmr_registers(1)(417)    <= not(local_tmr_voter(416));                                                                           
                tmr_registers(2)(417)    <= not(local_tmr_voter(416));                                                                           
 
                tmr_registers(0)(418)    <= not(local_tmr_voter(417));                                                                           
                tmr_registers(1)(418)    <= not(local_tmr_voter(417));                                                                           
                tmr_registers(2)(418)    <= not(local_tmr_voter(417));                                                                           
 
                tmr_registers(0)(419)    <= not(local_tmr_voter(418));                                                                           
                tmr_registers(1)(419)    <= not(local_tmr_voter(418));                                                                           
                tmr_registers(2)(419)    <= not(local_tmr_voter(418));                                                                           
 
                tmr_registers(0)(420)    <= not(local_tmr_voter(419));                                                                           
                tmr_registers(1)(420)    <= not(local_tmr_voter(419));                                                                           
                tmr_registers(2)(420)    <= not(local_tmr_voter(419));                                                                           
 
                tmr_registers(0)(421)    <= not(local_tmr_voter(420));                                                                           
                tmr_registers(1)(421)    <= not(local_tmr_voter(420));                                                                           
                tmr_registers(2)(421)    <= not(local_tmr_voter(420));                                                                           
 
                tmr_registers(0)(422)    <= not(local_tmr_voter(421));                                                                           
                tmr_registers(1)(422)    <= not(local_tmr_voter(421));                                                                           
                tmr_registers(2)(422)    <= not(local_tmr_voter(421));                                                                           
 
                tmr_registers(0)(423)    <= not(local_tmr_voter(422));                                                                           
                tmr_registers(1)(423)    <= not(local_tmr_voter(422));                                                                           
                tmr_registers(2)(423)    <= not(local_tmr_voter(422));                                                                           
 
                tmr_registers(0)(424)    <= not(local_tmr_voter(423));                                                                           
                tmr_registers(1)(424)    <= not(local_tmr_voter(423));                                                                           
                tmr_registers(2)(424)    <= not(local_tmr_voter(423));                                                                           
 
                tmr_registers(0)(425)    <= not(local_tmr_voter(424));                                                                           
                tmr_registers(1)(425)    <= not(local_tmr_voter(424));                                                                           
                tmr_registers(2)(425)    <= not(local_tmr_voter(424));                                                                           
 
                tmr_registers(0)(426)    <= not(local_tmr_voter(425));                                                                           
                tmr_registers(1)(426)    <= not(local_tmr_voter(425));                                                                           
                tmr_registers(2)(426)    <= not(local_tmr_voter(425));                                                                           
 
                tmr_registers(0)(427)    <= not(local_tmr_voter(426));                                                                           
                tmr_registers(1)(427)    <= not(local_tmr_voter(426));                                                                           
                tmr_registers(2)(427)    <= not(local_tmr_voter(426));                                                                           
 
                tmr_registers(0)(428)    <= not(local_tmr_voter(427));                                                                           
                tmr_registers(1)(428)    <= not(local_tmr_voter(427));                                                                           
                tmr_registers(2)(428)    <= not(local_tmr_voter(427));                                                                           
 
                tmr_registers(0)(429)    <= not(local_tmr_voter(428));                                                                           
                tmr_registers(1)(429)    <= not(local_tmr_voter(428));                                                                           
                tmr_registers(2)(429)    <= not(local_tmr_voter(428));                                                                           
 
                tmr_registers(0)(430)    <= not(local_tmr_voter(429));                                                                           
                tmr_registers(1)(430)    <= not(local_tmr_voter(429));                                                                           
                tmr_registers(2)(430)    <= not(local_tmr_voter(429));                                                                           
 
                tmr_registers(0)(431)    <= not(local_tmr_voter(430));                                                                           
                tmr_registers(1)(431)    <= not(local_tmr_voter(430));                                                                           
                tmr_registers(2)(431)    <= not(local_tmr_voter(430));                                                                           
 
                tmr_registers(0)(432)    <= not(local_tmr_voter(431));                                                                           
                tmr_registers(1)(432)    <= not(local_tmr_voter(431));                                                                           
                tmr_registers(2)(432)    <= not(local_tmr_voter(431));                                                                           
 
                tmr_registers(0)(433)    <= not(local_tmr_voter(432));                                                                           
                tmr_registers(1)(433)    <= not(local_tmr_voter(432));                                                                           
                tmr_registers(2)(433)    <= not(local_tmr_voter(432));                                                                           
 
                tmr_registers(0)(434)    <= not(local_tmr_voter(433));                                                                           
                tmr_registers(1)(434)    <= not(local_tmr_voter(433));                                                                           
                tmr_registers(2)(434)    <= not(local_tmr_voter(433));                                                                           
 
                tmr_registers(0)(435)    <= not(local_tmr_voter(434));                                                                           
                tmr_registers(1)(435)    <= not(local_tmr_voter(434));                                                                           
                tmr_registers(2)(435)    <= not(local_tmr_voter(434));                                                                           
 
                tmr_registers(0)(436)    <= not(local_tmr_voter(435));                                                                           
                tmr_registers(1)(436)    <= not(local_tmr_voter(435));                                                                           
                tmr_registers(2)(436)    <= not(local_tmr_voter(435));                                                                           
 
                tmr_registers(0)(437)    <= not(local_tmr_voter(436));                                                                           
                tmr_registers(1)(437)    <= not(local_tmr_voter(436));                                                                           
                tmr_registers(2)(437)    <= not(local_tmr_voter(436));                                                                           
 
                tmr_registers(0)(438)    <= not(local_tmr_voter(437));                                                                           
                tmr_registers(1)(438)    <= not(local_tmr_voter(437));                                                                           
                tmr_registers(2)(438)    <= not(local_tmr_voter(437));                                                                           
 
                tmr_registers(0)(439)    <= not(local_tmr_voter(438));                                                                           
                tmr_registers(1)(439)    <= not(local_tmr_voter(438));                                                                           
                tmr_registers(2)(439)    <= not(local_tmr_voter(438));                                                                           
 
                tmr_registers(0)(440)    <= not(local_tmr_voter(439));                                                                           
                tmr_registers(1)(440)    <= not(local_tmr_voter(439));                                                                           
                tmr_registers(2)(440)    <= not(local_tmr_voter(439));                                                                           
 
                tmr_registers(0)(441)    <= not(local_tmr_voter(440));                                                                           
                tmr_registers(1)(441)    <= not(local_tmr_voter(440));                                                                           
                tmr_registers(2)(441)    <= not(local_tmr_voter(440));                                                                           
 
                tmr_registers(0)(442)    <= not(local_tmr_voter(441));                                                                           
                tmr_registers(1)(442)    <= not(local_tmr_voter(441));                                                                           
                tmr_registers(2)(442)    <= not(local_tmr_voter(441));                                                                           
 
                tmr_registers(0)(443)    <= not(local_tmr_voter(442));                                                                           
                tmr_registers(1)(443)    <= not(local_tmr_voter(442));                                                                           
                tmr_registers(2)(443)    <= not(local_tmr_voter(442));                                                                           
 
                tmr_registers(0)(444)    <= not(local_tmr_voter(443));                                                                           
                tmr_registers(1)(444)    <= not(local_tmr_voter(443));                                                                           
                tmr_registers(2)(444)    <= not(local_tmr_voter(443));                                                                           
 
                tmr_registers(0)(445)    <= not(local_tmr_voter(444));                                                                           
                tmr_registers(1)(445)    <= not(local_tmr_voter(444));                                                                           
                tmr_registers(2)(445)    <= not(local_tmr_voter(444));                                                                           
 
                tmr_registers(0)(446)    <= not(local_tmr_voter(445));                                                                           
                tmr_registers(1)(446)    <= not(local_tmr_voter(445));                                                                           
                tmr_registers(2)(446)    <= not(local_tmr_voter(445));                                                                           
 
                tmr_registers(0)(447)    <= not(local_tmr_voter(446));                                                                           
                tmr_registers(1)(447)    <= not(local_tmr_voter(446));                                                                           
                tmr_registers(2)(447)    <= not(local_tmr_voter(446));                                                                           
 
                tmr_registers(0)(448)    <= not(local_tmr_voter(447));                                                                           
                tmr_registers(1)(448)    <= not(local_tmr_voter(447));                                                                           
                tmr_registers(2)(448)    <= not(local_tmr_voter(447));                                                                           
 
                tmr_registers(0)(449)    <= not(local_tmr_voter(448));                                                                           
                tmr_registers(1)(449)    <= not(local_tmr_voter(448));                                                                           
                tmr_registers(2)(449)    <= not(local_tmr_voter(448));                                                                           
 
                tmr_registers(0)(450)    <= not(local_tmr_voter(449));                                                                           
                tmr_registers(1)(450)    <= not(local_tmr_voter(449));                                                                           
                tmr_registers(2)(450)    <= not(local_tmr_voter(449));                                                                           
 
                tmr_registers(0)(451)    <= not(local_tmr_voter(450));                                                                           
                tmr_registers(1)(451)    <= not(local_tmr_voter(450));                                                                           
                tmr_registers(2)(451)    <= not(local_tmr_voter(450));                                                                           
 
                tmr_registers(0)(452)    <= not(local_tmr_voter(451));                                                                           
                tmr_registers(1)(452)    <= not(local_tmr_voter(451));                                                                           
                tmr_registers(2)(452)    <= not(local_tmr_voter(451));                                                                           
 
                tmr_registers(0)(453)    <= not(local_tmr_voter(452));                                                                           
                tmr_registers(1)(453)    <= not(local_tmr_voter(452));                                                                           
                tmr_registers(2)(453)    <= not(local_tmr_voter(452));                                                                           
 
                tmr_registers(0)(454)    <= not(local_tmr_voter(453));                                                                           
                tmr_registers(1)(454)    <= not(local_tmr_voter(453));                                                                           
                tmr_registers(2)(454)    <= not(local_tmr_voter(453));                                                                           
 
                tmr_registers(0)(455)    <= not(local_tmr_voter(454));                                                                           
                tmr_registers(1)(455)    <= not(local_tmr_voter(454));                                                                           
                tmr_registers(2)(455)    <= not(local_tmr_voter(454));                                                                           
 
                tmr_registers(0)(456)    <= not(local_tmr_voter(455));                                                                           
                tmr_registers(1)(456)    <= not(local_tmr_voter(455));                                                                           
                tmr_registers(2)(456)    <= not(local_tmr_voter(455));                                                                           
 
                tmr_registers(0)(457)    <= not(local_tmr_voter(456));                                                                           
                tmr_registers(1)(457)    <= not(local_tmr_voter(456));                                                                           
                tmr_registers(2)(457)    <= not(local_tmr_voter(456));                                                                           
 
                tmr_registers(0)(458)    <= not(local_tmr_voter(457));                                                                           
                tmr_registers(1)(458)    <= not(local_tmr_voter(457));                                                                           
                tmr_registers(2)(458)    <= not(local_tmr_voter(457));                                                                           
 
                tmr_registers(0)(459)    <= not(local_tmr_voter(458));                                                                           
                tmr_registers(1)(459)    <= not(local_tmr_voter(458));                                                                           
                tmr_registers(2)(459)    <= not(local_tmr_voter(458));                                                                           
 
                tmr_registers(0)(460)    <= not(local_tmr_voter(459));                                                                           
                tmr_registers(1)(460)    <= not(local_tmr_voter(459));                                                                           
                tmr_registers(2)(460)    <= not(local_tmr_voter(459));                                                                           
 
                tmr_registers(0)(461)    <= not(local_tmr_voter(460));                                                                           
                tmr_registers(1)(461)    <= not(local_tmr_voter(460));                                                                           
                tmr_registers(2)(461)    <= not(local_tmr_voter(460));                                                                           
 
                tmr_registers(0)(462)    <= not(local_tmr_voter(461));                                                                           
                tmr_registers(1)(462)    <= not(local_tmr_voter(461));                                                                           
                tmr_registers(2)(462)    <= not(local_tmr_voter(461));                                                                           
 
                tmr_registers(0)(463)    <= not(local_tmr_voter(462));                                                                           
                tmr_registers(1)(463)    <= not(local_tmr_voter(462));                                                                           
                tmr_registers(2)(463)    <= not(local_tmr_voter(462));                                                                           
 
                tmr_registers(0)(464)    <= not(local_tmr_voter(463));                                                                           
                tmr_registers(1)(464)    <= not(local_tmr_voter(463));                                                                           
                tmr_registers(2)(464)    <= not(local_tmr_voter(463));                                                                           
 
                tmr_registers(0)(465)    <= not(local_tmr_voter(464));                                                                           
                tmr_registers(1)(465)    <= not(local_tmr_voter(464));                                                                           
                tmr_registers(2)(465)    <= not(local_tmr_voter(464));                                                                           
 
                tmr_registers(0)(466)    <= not(local_tmr_voter(465));                                                                           
                tmr_registers(1)(466)    <= not(local_tmr_voter(465));                                                                           
                tmr_registers(2)(466)    <= not(local_tmr_voter(465));                                                                           
 
                tmr_registers(0)(467)    <= not(local_tmr_voter(466));                                                                           
                tmr_registers(1)(467)    <= not(local_tmr_voter(466));                                                                           
                tmr_registers(2)(467)    <= not(local_tmr_voter(466));                                                                           
 
                tmr_registers(0)(468)    <= not(local_tmr_voter(467));                                                                           
                tmr_registers(1)(468)    <= not(local_tmr_voter(467));                                                                           
                tmr_registers(2)(468)    <= not(local_tmr_voter(467));                                                                           
 
                tmr_registers(0)(469)    <= not(local_tmr_voter(468));                                                                           
                tmr_registers(1)(469)    <= not(local_tmr_voter(468));                                                                           
                tmr_registers(2)(469)    <= not(local_tmr_voter(468));                                                                           
 
                tmr_registers(0)(470)    <= not(local_tmr_voter(469));                                                                           
                tmr_registers(1)(470)    <= not(local_tmr_voter(469));                                                                           
                tmr_registers(2)(470)    <= not(local_tmr_voter(469));                                                                           
 
                tmr_registers(0)(471)    <= not(local_tmr_voter(470));                                                                           
                tmr_registers(1)(471)    <= not(local_tmr_voter(470));                                                                           
                tmr_registers(2)(471)    <= not(local_tmr_voter(470));                                                                           
 
                tmr_registers(0)(472)    <= not(local_tmr_voter(471));                                                                           
                tmr_registers(1)(472)    <= not(local_tmr_voter(471));                                                                           
                tmr_registers(2)(472)    <= not(local_tmr_voter(471));                                                                           
 
                tmr_registers(0)(473)    <= not(local_tmr_voter(472));                                                                           
                tmr_registers(1)(473)    <= not(local_tmr_voter(472));                                                                           
                tmr_registers(2)(473)    <= not(local_tmr_voter(472));                                                                           
 
                tmr_registers(0)(474)    <= not(local_tmr_voter(473));                                                                           
                tmr_registers(1)(474)    <= not(local_tmr_voter(473));                                                                           
                tmr_registers(2)(474)    <= not(local_tmr_voter(473));                                                                           
 
                tmr_registers(0)(475)    <= not(local_tmr_voter(474));                                                                           
                tmr_registers(1)(475)    <= not(local_tmr_voter(474));                                                                           
                tmr_registers(2)(475)    <= not(local_tmr_voter(474));                                                                           
 
                tmr_registers(0)(476)    <= not(local_tmr_voter(475));                                                                           
                tmr_registers(1)(476)    <= not(local_tmr_voter(475));                                                                           
                tmr_registers(2)(476)    <= not(local_tmr_voter(475));                                                                           
 
                tmr_registers(0)(477)    <= not(local_tmr_voter(476));                                                                           
                tmr_registers(1)(477)    <= not(local_tmr_voter(476));                                                                           
                tmr_registers(2)(477)    <= not(local_tmr_voter(476));                                                                           
 
                tmr_registers(0)(478)    <= not(local_tmr_voter(477));                                                                           
                tmr_registers(1)(478)    <= not(local_tmr_voter(477));                                                                           
                tmr_registers(2)(478)    <= not(local_tmr_voter(477));                                                                           
 
                tmr_registers(0)(479)    <= not(local_tmr_voter(478));                                                                           
                tmr_registers(1)(479)    <= not(local_tmr_voter(478));                                                                           
                tmr_registers(2)(479)    <= not(local_tmr_voter(478));                                                                           
 
                tmr_registers(0)(480)    <= not(local_tmr_voter(479));                                                                           
                tmr_registers(1)(480)    <= not(local_tmr_voter(479));                                                                           
                tmr_registers(2)(480)    <= not(local_tmr_voter(479));                                                                           
 
                tmr_registers(0)(481)    <= not(local_tmr_voter(480));                                                                           
                tmr_registers(1)(481)    <= not(local_tmr_voter(480));                                                                           
                tmr_registers(2)(481)    <= not(local_tmr_voter(480));                                                                           
 
                tmr_registers(0)(482)    <= not(local_tmr_voter(481));                                                                           
                tmr_registers(1)(482)    <= not(local_tmr_voter(481));                                                                           
                tmr_registers(2)(482)    <= not(local_tmr_voter(481));                                                                           
 
                tmr_registers(0)(483)    <= not(local_tmr_voter(482));                                                                           
                tmr_registers(1)(483)    <= not(local_tmr_voter(482));                                                                           
                tmr_registers(2)(483)    <= not(local_tmr_voter(482));                                                                           
 
                tmr_registers(0)(484)    <= not(local_tmr_voter(483));                                                                           
                tmr_registers(1)(484)    <= not(local_tmr_voter(483));                                                                           
                tmr_registers(2)(484)    <= not(local_tmr_voter(483));                                                                           
 
                tmr_registers(0)(485)    <= not(local_tmr_voter(484));                                                                           
                tmr_registers(1)(485)    <= not(local_tmr_voter(484));                                                                           
                tmr_registers(2)(485)    <= not(local_tmr_voter(484));                                                                           
 
                tmr_registers(0)(486)    <= not(local_tmr_voter(485));                                                                           
                tmr_registers(1)(486)    <= not(local_tmr_voter(485));                                                                           
                tmr_registers(2)(486)    <= not(local_tmr_voter(485));                                                                           
 
                tmr_registers(0)(487)    <= not(local_tmr_voter(486));                                                                           
                tmr_registers(1)(487)    <= not(local_tmr_voter(486));                                                                           
                tmr_registers(2)(487)    <= not(local_tmr_voter(486));                                                                           
 
                tmr_registers(0)(488)    <= not(local_tmr_voter(487));                                                                           
                tmr_registers(1)(488)    <= not(local_tmr_voter(487));                                                                           
                tmr_registers(2)(488)    <= not(local_tmr_voter(487));                                                                           
 
                tmr_registers(0)(489)    <= not(local_tmr_voter(488));                                                                           
                tmr_registers(1)(489)    <= not(local_tmr_voter(488));                                                                           
                tmr_registers(2)(489)    <= not(local_tmr_voter(488));                                                                           
 
                tmr_registers(0)(490)    <= not(local_tmr_voter(489));                                                                           
                tmr_registers(1)(490)    <= not(local_tmr_voter(489));                                                                           
                tmr_registers(2)(490)    <= not(local_tmr_voter(489));                                                                           
 
                tmr_registers(0)(491)    <= not(local_tmr_voter(490));                                                                           
                tmr_registers(1)(491)    <= not(local_tmr_voter(490));                                                                           
                tmr_registers(2)(491)    <= not(local_tmr_voter(490));                                                                           
 
                tmr_registers(0)(492)    <= not(local_tmr_voter(491));                                                                           
                tmr_registers(1)(492)    <= not(local_tmr_voter(491));                                                                           
                tmr_registers(2)(492)    <= not(local_tmr_voter(491));                                                                           
 
                tmr_registers(0)(493)    <= not(local_tmr_voter(492));                                                                           
                tmr_registers(1)(493)    <= not(local_tmr_voter(492));                                                                           
                tmr_registers(2)(493)    <= not(local_tmr_voter(492));                                                                           
 
                tmr_registers(0)(494)    <= not(local_tmr_voter(493));                                                                           
                tmr_registers(1)(494)    <= not(local_tmr_voter(493));                                                                           
                tmr_registers(2)(494)    <= not(local_tmr_voter(493));                                                                           
 
                tmr_registers(0)(495)    <= not(local_tmr_voter(494));                                                                           
                tmr_registers(1)(495)    <= not(local_tmr_voter(494));                                                                           
                tmr_registers(2)(495)    <= not(local_tmr_voter(494));                                                                           
 
                tmr_registers(0)(496)    <= not(local_tmr_voter(495));                                                                           
                tmr_registers(1)(496)    <= not(local_tmr_voter(495));                                                                           
                tmr_registers(2)(496)    <= not(local_tmr_voter(495));                                                                           
 
                tmr_registers(0)(497)    <= not(local_tmr_voter(496));                                                                           
                tmr_registers(1)(497)    <= not(local_tmr_voter(496));                                                                           
                tmr_registers(2)(497)    <= not(local_tmr_voter(496));                                                                           
 
                tmr_registers(0)(498)    <= not(local_tmr_voter(497));                                                                           
                tmr_registers(1)(498)    <= not(local_tmr_voter(497));                                                                           
                tmr_registers(2)(498)    <= not(local_tmr_voter(497));                                                                           
 
                tmr_registers(0)(499)    <= not(local_tmr_voter(498));                                                                           
                tmr_registers(1)(499)    <= not(local_tmr_voter(498));                                                                           
                tmr_registers(2)(499)    <= not(local_tmr_voter(498));                                                                           
 
                tmr_registers(0)(500)    <= not(local_tmr_voter(499));                                                                           
                tmr_registers(1)(500)    <= not(local_tmr_voter(499));                                                                           
                tmr_registers(2)(500)    <= not(local_tmr_voter(499));                                                                           
 
                tmr_registers(0)(501)    <= not(local_tmr_voter(500));                                                                           
                tmr_registers(1)(501)    <= not(local_tmr_voter(500));                                                                           
                tmr_registers(2)(501)    <= not(local_tmr_voter(500));                                                                           
 
                tmr_registers(0)(502)    <= not(local_tmr_voter(501));                                                                           
                tmr_registers(1)(502)    <= not(local_tmr_voter(501));                                                                           
                tmr_registers(2)(502)    <= not(local_tmr_voter(501));                                                                           
 
                tmr_registers(0)(503)    <= not(local_tmr_voter(502));                                                                           
                tmr_registers(1)(503)    <= not(local_tmr_voter(502));                                                                           
                tmr_registers(2)(503)    <= not(local_tmr_voter(502));                                                                           
 
                tmr_registers(0)(504)    <= not(local_tmr_voter(503));                                                                           
                tmr_registers(1)(504)    <= not(local_tmr_voter(503));                                                                           
                tmr_registers(2)(504)    <= not(local_tmr_voter(503));                                                                           
 
                tmr_registers(0)(505)    <= not(local_tmr_voter(504));                                                                           
                tmr_registers(1)(505)    <= not(local_tmr_voter(504));                                                                           
                tmr_registers(2)(505)    <= not(local_tmr_voter(504));                                                                           
 
                tmr_registers(0)(506)    <= not(local_tmr_voter(505));                                                                           
                tmr_registers(1)(506)    <= not(local_tmr_voter(505));                                                                           
                tmr_registers(2)(506)    <= not(local_tmr_voter(505));                                                                           
 
                tmr_registers(0)(507)    <= not(local_tmr_voter(506));                                                                           
                tmr_registers(1)(507)    <= not(local_tmr_voter(506));                                                                           
                tmr_registers(2)(507)    <= not(local_tmr_voter(506));                                                                           
 
                tmr_registers(0)(508)    <= not(local_tmr_voter(507));                                                                           
                tmr_registers(1)(508)    <= not(local_tmr_voter(507));                                                                           
                tmr_registers(2)(508)    <= not(local_tmr_voter(507));                                                                           
 
                tmr_registers(0)(509)    <= not(local_tmr_voter(508));                                                                           
                tmr_registers(1)(509)    <= not(local_tmr_voter(508));                                                                           
                tmr_registers(2)(509)    <= not(local_tmr_voter(508));                                                                           
 
                tmr_registers(0)(510)    <= not(local_tmr_voter(509));                                                                           
                tmr_registers(1)(510)    <= not(local_tmr_voter(509));                                                                           
                tmr_registers(2)(510)    <= not(local_tmr_voter(509));                                                                           
 
                tmr_registers(0)(511)    <= not(local_tmr_voter(510));                                                                           
                tmr_registers(1)(511)    <= not(local_tmr_voter(510));                                                                           
                tmr_registers(2)(511)    <= not(local_tmr_voter(510));                                                                           
 
                tmr_registers(0)(512)    <= not(local_tmr_voter(511));                                                                           
                tmr_registers(1)(512)    <= not(local_tmr_voter(511));                                                                           
                tmr_registers(2)(512)    <= not(local_tmr_voter(511));                                                                           
 
                tmr_registers(0)(513)    <= not(local_tmr_voter(512));                                                                           
                tmr_registers(1)(513)    <= not(local_tmr_voter(512));                                                                           
                tmr_registers(2)(513)    <= not(local_tmr_voter(512));                                                                           
 
                tmr_registers(0)(514)    <= not(local_tmr_voter(513));                                                                           
                tmr_registers(1)(514)    <= not(local_tmr_voter(513));                                                                           
                tmr_registers(2)(514)    <= not(local_tmr_voter(513));                                                                           
 
                tmr_registers(0)(515)    <= not(local_tmr_voter(514));                                                                           
                tmr_registers(1)(515)    <= not(local_tmr_voter(514));                                                                           
                tmr_registers(2)(515)    <= not(local_tmr_voter(514));                                                                           
 
                tmr_registers(0)(516)    <= not(local_tmr_voter(515));                                                                           
                tmr_registers(1)(516)    <= not(local_tmr_voter(515));                                                                           
                tmr_registers(2)(516)    <= not(local_tmr_voter(515));                                                                           
 
                tmr_registers(0)(517)    <= not(local_tmr_voter(516));                                                                           
                tmr_registers(1)(517)    <= not(local_tmr_voter(516));                                                                           
                tmr_registers(2)(517)    <= not(local_tmr_voter(516));                                                                           
 
                tmr_registers(0)(518)    <= not(local_tmr_voter(517));                                                                           
                tmr_registers(1)(518)    <= not(local_tmr_voter(517));                                                                           
                tmr_registers(2)(518)    <= not(local_tmr_voter(517));                                                                           
 
                tmr_registers(0)(519)    <= not(local_tmr_voter(518));                                                                           
                tmr_registers(1)(519)    <= not(local_tmr_voter(518));                                                                           
                tmr_registers(2)(519)    <= not(local_tmr_voter(518));                                                                           
 
                tmr_registers(0)(520)    <= not(local_tmr_voter(519));                                                                           
                tmr_registers(1)(520)    <= not(local_tmr_voter(519));                                                                           
                tmr_registers(2)(520)    <= not(local_tmr_voter(519));                                                                           
 
                tmr_registers(0)(521)    <= not(local_tmr_voter(520));                                                                           
                tmr_registers(1)(521)    <= not(local_tmr_voter(520));                                                                           
                tmr_registers(2)(521)    <= not(local_tmr_voter(520));                                                                           
 
                tmr_registers(0)(522)    <= not(local_tmr_voter(521));                                                                           
                tmr_registers(1)(522)    <= not(local_tmr_voter(521));                                                                           
                tmr_registers(2)(522)    <= not(local_tmr_voter(521));                                                                           
 
                tmr_registers(0)(523)    <= not(local_tmr_voter(522));                                                                           
                tmr_registers(1)(523)    <= not(local_tmr_voter(522));                                                                           
                tmr_registers(2)(523)    <= not(local_tmr_voter(522));                                                                           
 
                tmr_registers(0)(524)    <= not(local_tmr_voter(523));                                                                           
                tmr_registers(1)(524)    <= not(local_tmr_voter(523));                                                                           
                tmr_registers(2)(524)    <= not(local_tmr_voter(523));                                                                           
 
                tmr_registers(0)(525)    <= not(local_tmr_voter(524));                                                                           
                tmr_registers(1)(525)    <= not(local_tmr_voter(524));                                                                           
                tmr_registers(2)(525)    <= not(local_tmr_voter(524));                                                                           
 
                tmr_registers(0)(526)    <= not(local_tmr_voter(525));                                                                           
                tmr_registers(1)(526)    <= not(local_tmr_voter(525));                                                                           
                tmr_registers(2)(526)    <= not(local_tmr_voter(525));                                                                           
 
                tmr_registers(0)(527)    <= not(local_tmr_voter(526));                                                                           
                tmr_registers(1)(527)    <= not(local_tmr_voter(526));                                                                           
                tmr_registers(2)(527)    <= not(local_tmr_voter(526));                                                                           
 
                tmr_registers(0)(528)    <= not(local_tmr_voter(527));                                                                           
                tmr_registers(1)(528)    <= not(local_tmr_voter(527));                                                                           
                tmr_registers(2)(528)    <= not(local_tmr_voter(527));                                                                           
 
                tmr_registers(0)(529)    <= not(local_tmr_voter(528));                                                                           
                tmr_registers(1)(529)    <= not(local_tmr_voter(528));                                                                           
                tmr_registers(2)(529)    <= not(local_tmr_voter(528));                                                                           
 
                tmr_registers(0)(530)    <= not(local_tmr_voter(529));                                                                           
                tmr_registers(1)(530)    <= not(local_tmr_voter(529));                                                                           
                tmr_registers(2)(530)    <= not(local_tmr_voter(529));                                                                           
 
                tmr_registers(0)(531)    <= not(local_tmr_voter(530));                                                                           
                tmr_registers(1)(531)    <= not(local_tmr_voter(530));                                                                           
                tmr_registers(2)(531)    <= not(local_tmr_voter(530));                                                                           
 
                tmr_registers(0)(532)    <= not(local_tmr_voter(531));                                                                           
                tmr_registers(1)(532)    <= not(local_tmr_voter(531));                                                                           
                tmr_registers(2)(532)    <= not(local_tmr_voter(531));                                                                           
 
                tmr_registers(0)(533)    <= not(local_tmr_voter(532));                                                                           
                tmr_registers(1)(533)    <= not(local_tmr_voter(532));                                                                           
                tmr_registers(2)(533)    <= not(local_tmr_voter(532));                                                                           
 
                tmr_registers(0)(534)    <= not(local_tmr_voter(533));                                                                           
                tmr_registers(1)(534)    <= not(local_tmr_voter(533));                                                                           
                tmr_registers(2)(534)    <= not(local_tmr_voter(533));                                                                           
 
                tmr_registers(0)(535)    <= not(local_tmr_voter(534));                                                                           
                tmr_registers(1)(535)    <= not(local_tmr_voter(534));                                                                           
                tmr_registers(2)(535)    <= not(local_tmr_voter(534));                                                                           
 
                tmr_registers(0)(536)    <= not(local_tmr_voter(535));                                                                           
                tmr_registers(1)(536)    <= not(local_tmr_voter(535));                                                                           
                tmr_registers(2)(536)    <= not(local_tmr_voter(535));                                                                           
 
                tmr_registers(0)(537)    <= not(local_tmr_voter(536));                                                                           
                tmr_registers(1)(537)    <= not(local_tmr_voter(536));                                                                           
                tmr_registers(2)(537)    <= not(local_tmr_voter(536));                                                                           
 
                tmr_registers(0)(538)    <= not(local_tmr_voter(537));                                                                           
                tmr_registers(1)(538)    <= not(local_tmr_voter(537));                                                                           
                tmr_registers(2)(538)    <= not(local_tmr_voter(537));                                                                           
 
                tmr_registers(0)(539)    <= not(local_tmr_voter(538));                                                                           
                tmr_registers(1)(539)    <= not(local_tmr_voter(538));                                                                           
                tmr_registers(2)(539)    <= not(local_tmr_voter(538));                                                                           
 
                tmr_registers(0)(540)    <= not(local_tmr_voter(539));                                                                           
                tmr_registers(1)(540)    <= not(local_tmr_voter(539));                                                                           
                tmr_registers(2)(540)    <= not(local_tmr_voter(539));                                                                           
 
                tmr_registers(0)(541)    <= not(local_tmr_voter(540));                                                                           
                tmr_registers(1)(541)    <= not(local_tmr_voter(540));                                                                           
                tmr_registers(2)(541)    <= not(local_tmr_voter(540));                                                                           
 
                tmr_registers(0)(542)    <= not(local_tmr_voter(541));                                                                           
                tmr_registers(1)(542)    <= not(local_tmr_voter(541));                                                                           
                tmr_registers(2)(542)    <= not(local_tmr_voter(541));                                                                           
 
                tmr_registers(0)(543)    <= not(local_tmr_voter(542));                                                                           
                tmr_registers(1)(543)    <= not(local_tmr_voter(542));                                                                           
                tmr_registers(2)(543)    <= not(local_tmr_voter(542));                                                                           
 
                tmr_registers(0)(544)    <= not(local_tmr_voter(543));                                                                           
                tmr_registers(1)(544)    <= not(local_tmr_voter(543));                                                                           
                tmr_registers(2)(544)    <= not(local_tmr_voter(543));                                                                           
 
                tmr_registers(0)(545)    <= not(local_tmr_voter(544));                                                                           
                tmr_registers(1)(545)    <= not(local_tmr_voter(544));                                                                           
                tmr_registers(2)(545)    <= not(local_tmr_voter(544));                                                                           
 
                tmr_registers(0)(546)    <= not(local_tmr_voter(545));                                                                           
                tmr_registers(1)(546)    <= not(local_tmr_voter(545));                                                                           
                tmr_registers(2)(546)    <= not(local_tmr_voter(545));                                                                           
 
                tmr_registers(0)(547)    <= not(local_tmr_voter(546));                                                                           
                tmr_registers(1)(547)    <= not(local_tmr_voter(546));                                                                           
                tmr_registers(2)(547)    <= not(local_tmr_voter(546));                                                                           
 
                tmr_registers(0)(548)    <= not(local_tmr_voter(547));                                                                           
                tmr_registers(1)(548)    <= not(local_tmr_voter(547));                                                                           
                tmr_registers(2)(548)    <= not(local_tmr_voter(547));                                                                           
 
                tmr_registers(0)(549)    <= not(local_tmr_voter(548));                                                                           
                tmr_registers(1)(549)    <= not(local_tmr_voter(548));                                                                           
                tmr_registers(2)(549)    <= not(local_tmr_voter(548));                                                                           
 
                tmr_registers(0)(550)    <= not(local_tmr_voter(549));                                                                           
                tmr_registers(1)(550)    <= not(local_tmr_voter(549));                                                                           
                tmr_registers(2)(550)    <= not(local_tmr_voter(549));                                                                           
 
                tmr_registers(0)(551)    <= not(local_tmr_voter(550));                                                                           
                tmr_registers(1)(551)    <= not(local_tmr_voter(550));                                                                           
                tmr_registers(2)(551)    <= not(local_tmr_voter(550));                                                                           
 
                tmr_registers(0)(552)    <= not(local_tmr_voter(551));                                                                           
                tmr_registers(1)(552)    <= not(local_tmr_voter(551));                                                                           
                tmr_registers(2)(552)    <= not(local_tmr_voter(551));                                                                           
 
                tmr_registers(0)(553)    <= not(local_tmr_voter(552));                                                                           
                tmr_registers(1)(553)    <= not(local_tmr_voter(552));                                                                           
                tmr_registers(2)(553)    <= not(local_tmr_voter(552));                                                                           
 
                tmr_registers(0)(554)    <= not(local_tmr_voter(553));                                                                           
                tmr_registers(1)(554)    <= not(local_tmr_voter(553));                                                                           
                tmr_registers(2)(554)    <= not(local_tmr_voter(553));                                                                           
 
                tmr_registers(0)(555)    <= not(local_tmr_voter(554));                                                                           
                tmr_registers(1)(555)    <= not(local_tmr_voter(554));                                                                           
                tmr_registers(2)(555)    <= not(local_tmr_voter(554));                                                                           
 
                tmr_registers(0)(556)    <= not(local_tmr_voter(555));                                                                           
                tmr_registers(1)(556)    <= not(local_tmr_voter(555));                                                                           
                tmr_registers(2)(556)    <= not(local_tmr_voter(555));                                                                           
 
                tmr_registers(0)(557)    <= not(local_tmr_voter(556));                                                                           
                tmr_registers(1)(557)    <= not(local_tmr_voter(556));                                                                           
                tmr_registers(2)(557)    <= not(local_tmr_voter(556));                                                                           
 
                tmr_registers(0)(558)    <= not(local_tmr_voter(557));                                                                           
                tmr_registers(1)(558)    <= not(local_tmr_voter(557));                                                                           
                tmr_registers(2)(558)    <= not(local_tmr_voter(557));                                                                           
 
                tmr_registers(0)(559)    <= not(local_tmr_voter(558));                                                                           
                tmr_registers(1)(559)    <= not(local_tmr_voter(558));                                                                           
                tmr_registers(2)(559)    <= not(local_tmr_voter(558));                                                                           
 
                tmr_registers(0)(560)    <= not(local_tmr_voter(559));                                                                           
                tmr_registers(1)(560)    <= not(local_tmr_voter(559));                                                                           
                tmr_registers(2)(560)    <= not(local_tmr_voter(559));                                                                           
 
                tmr_registers(0)(561)    <= not(local_tmr_voter(560));                                                                           
                tmr_registers(1)(561)    <= not(local_tmr_voter(560));                                                                           
                tmr_registers(2)(561)    <= not(local_tmr_voter(560));                                                                           
 
                tmr_registers(0)(562)    <= not(local_tmr_voter(561));                                                                           
                tmr_registers(1)(562)    <= not(local_tmr_voter(561));                                                                           
                tmr_registers(2)(562)    <= not(local_tmr_voter(561));                                                                           
 
                tmr_registers(0)(563)    <= not(local_tmr_voter(562));                                                                           
                tmr_registers(1)(563)    <= not(local_tmr_voter(562));                                                                           
                tmr_registers(2)(563)    <= not(local_tmr_voter(562));                                                                           
 
                tmr_registers(0)(564)    <= not(local_tmr_voter(563));                                                                           
                tmr_registers(1)(564)    <= not(local_tmr_voter(563));                                                                           
                tmr_registers(2)(564)    <= not(local_tmr_voter(563));                                                                           
 
                tmr_registers(0)(565)    <= not(local_tmr_voter(564));                                                                           
                tmr_registers(1)(565)    <= not(local_tmr_voter(564));                                                                           
                tmr_registers(2)(565)    <= not(local_tmr_voter(564));                                                                           
 
                tmr_registers(0)(566)    <= not(local_tmr_voter(565));                                                                           
                tmr_registers(1)(566)    <= not(local_tmr_voter(565));                                                                           
                tmr_registers(2)(566)    <= not(local_tmr_voter(565));                                                                           
 
                tmr_registers(0)(567)    <= not(local_tmr_voter(566));                                                                           
                tmr_registers(1)(567)    <= not(local_tmr_voter(566));                                                                           
                tmr_registers(2)(567)    <= not(local_tmr_voter(566));                                                                           
 
                tmr_registers(0)(568)    <= not(local_tmr_voter(567));                                                                           
                tmr_registers(1)(568)    <= not(local_tmr_voter(567));                                                                           
                tmr_registers(2)(568)    <= not(local_tmr_voter(567));                                                                           
 
                tmr_registers(0)(569)    <= not(local_tmr_voter(568));                                                                           
                tmr_registers(1)(569)    <= not(local_tmr_voter(568));                                                                           
                tmr_registers(2)(569)    <= not(local_tmr_voter(568));                                                                           
 
                tmr_registers(0)(570)    <= not(local_tmr_voter(569));                                                                           
                tmr_registers(1)(570)    <= not(local_tmr_voter(569));                                                                           
                tmr_registers(2)(570)    <= not(local_tmr_voter(569));                                                                           
 
                tmr_registers(0)(571)    <= not(local_tmr_voter(570));                                                                           
                tmr_registers(1)(571)    <= not(local_tmr_voter(570));                                                                           
                tmr_registers(2)(571)    <= not(local_tmr_voter(570));                                                                           
 
                tmr_registers(0)(572)    <= not(local_tmr_voter(571));                                                                           
                tmr_registers(1)(572)    <= not(local_tmr_voter(571));                                                                           
                tmr_registers(2)(572)    <= not(local_tmr_voter(571));                                                                           
 
                tmr_registers(0)(573)    <= not(local_tmr_voter(572));                                                                           
                tmr_registers(1)(573)    <= not(local_tmr_voter(572));                                                                           
                tmr_registers(2)(573)    <= not(local_tmr_voter(572));                                                                           
 
                tmr_registers(0)(574)    <= not(local_tmr_voter(573));                                                                           
                tmr_registers(1)(574)    <= not(local_tmr_voter(573));                                                                           
                tmr_registers(2)(574)    <= not(local_tmr_voter(573));                                                                           
 
                tmr_registers(0)(575)    <= not(local_tmr_voter(574));                                                                           
                tmr_registers(1)(575)    <= not(local_tmr_voter(574));                                                                           
                tmr_registers(2)(575)    <= not(local_tmr_voter(574));                                                                           
 
                tmr_registers(0)(576)    <= not(local_tmr_voter(575));                                                                           
                tmr_registers(1)(576)    <= not(local_tmr_voter(575));                                                                           
                tmr_registers(2)(576)    <= not(local_tmr_voter(575));                                                                           
 
                tmr_registers(0)(577)    <= not(local_tmr_voter(576));                                                                           
                tmr_registers(1)(577)    <= not(local_tmr_voter(576));                                                                           
                tmr_registers(2)(577)    <= not(local_tmr_voter(576));                                                                           
 
                tmr_registers(0)(578)    <= not(local_tmr_voter(577));                                                                           
                tmr_registers(1)(578)    <= not(local_tmr_voter(577));                                                                           
                tmr_registers(2)(578)    <= not(local_tmr_voter(577));                                                                           
 
                tmr_registers(0)(579)    <= not(local_tmr_voter(578));                                                                           
                tmr_registers(1)(579)    <= not(local_tmr_voter(578));                                                                           
                tmr_registers(2)(579)    <= not(local_tmr_voter(578));                                                                           
 
                tmr_registers(0)(580)    <= not(local_tmr_voter(579));                                                                           
                tmr_registers(1)(580)    <= not(local_tmr_voter(579));                                                                           
                tmr_registers(2)(580)    <= not(local_tmr_voter(579));                                                                           
 
                tmr_registers(0)(581)    <= not(local_tmr_voter(580));                                                                           
                tmr_registers(1)(581)    <= not(local_tmr_voter(580));                                                                           
                tmr_registers(2)(581)    <= not(local_tmr_voter(580));                                                                           
 
                tmr_registers(0)(582)    <= not(local_tmr_voter(581));                                                                           
                tmr_registers(1)(582)    <= not(local_tmr_voter(581));                                                                           
                tmr_registers(2)(582)    <= not(local_tmr_voter(581));                                                                           
 
                tmr_registers(0)(583)    <= not(local_tmr_voter(582));                                                                           
                tmr_registers(1)(583)    <= not(local_tmr_voter(582));                                                                           
                tmr_registers(2)(583)    <= not(local_tmr_voter(582));                                                                           
 
                tmr_registers(0)(584)    <= not(local_tmr_voter(583));                                                                           
                tmr_registers(1)(584)    <= not(local_tmr_voter(583));                                                                           
                tmr_registers(2)(584)    <= not(local_tmr_voter(583));                                                                           
 
                tmr_registers(0)(585)    <= not(local_tmr_voter(584));                                                                           
                tmr_registers(1)(585)    <= not(local_tmr_voter(584));                                                                           
                tmr_registers(2)(585)    <= not(local_tmr_voter(584));                                                                           
 
                tmr_registers(0)(586)    <= not(local_tmr_voter(585));                                                                           
                tmr_registers(1)(586)    <= not(local_tmr_voter(585));                                                                           
                tmr_registers(2)(586)    <= not(local_tmr_voter(585));                                                                           
 
                tmr_registers(0)(587)    <= not(local_tmr_voter(586));                                                                           
                tmr_registers(1)(587)    <= not(local_tmr_voter(586));                                                                           
                tmr_registers(2)(587)    <= not(local_tmr_voter(586));                                                                           
 
                tmr_registers(0)(588)    <= not(local_tmr_voter(587));                                                                           
                tmr_registers(1)(588)    <= not(local_tmr_voter(587));                                                                           
                tmr_registers(2)(588)    <= not(local_tmr_voter(587));                                                                           
 
                tmr_registers(0)(589)    <= not(local_tmr_voter(588));                                                                           
                tmr_registers(1)(589)    <= not(local_tmr_voter(588));                                                                           
                tmr_registers(2)(589)    <= not(local_tmr_voter(588));                                                                           
 
                tmr_registers(0)(590)    <= not(local_tmr_voter(589));                                                                           
                tmr_registers(1)(590)    <= not(local_tmr_voter(589));                                                                           
                tmr_registers(2)(590)    <= not(local_tmr_voter(589));                                                                           
 
                tmr_registers(0)(591)    <= not(local_tmr_voter(590));                                                                           
                tmr_registers(1)(591)    <= not(local_tmr_voter(590));                                                                           
                tmr_registers(2)(591)    <= not(local_tmr_voter(590));                                                                           
 
                tmr_registers(0)(592)    <= not(local_tmr_voter(591));                                                                           
                tmr_registers(1)(592)    <= not(local_tmr_voter(591));                                                                           
                tmr_registers(2)(592)    <= not(local_tmr_voter(591));                                                                           
 
                tmr_registers(0)(593)    <= not(local_tmr_voter(592));                                                                           
                tmr_registers(1)(593)    <= not(local_tmr_voter(592));                                                                           
                tmr_registers(2)(593)    <= not(local_tmr_voter(592));                                                                           
 
                tmr_registers(0)(594)    <= not(local_tmr_voter(593));                                                                           
                tmr_registers(1)(594)    <= not(local_tmr_voter(593));                                                                           
                tmr_registers(2)(594)    <= not(local_tmr_voter(593));                                                                           
 
                tmr_registers(0)(595)    <= not(local_tmr_voter(594));                                                                           
                tmr_registers(1)(595)    <= not(local_tmr_voter(594));                                                                           
                tmr_registers(2)(595)    <= not(local_tmr_voter(594));                                                                           
 
                tmr_registers(0)(596)    <= not(local_tmr_voter(595));                                                                           
                tmr_registers(1)(596)    <= not(local_tmr_voter(595));                                                                           
                tmr_registers(2)(596)    <= not(local_tmr_voter(595));                                                                           
 
                tmr_registers(0)(597)    <= not(local_tmr_voter(596));                                                                           
                tmr_registers(1)(597)    <= not(local_tmr_voter(596));                                                                           
                tmr_registers(2)(597)    <= not(local_tmr_voter(596));                                                                           
 
                tmr_registers(0)(598)    <= not(local_tmr_voter(597));                                                                           
                tmr_registers(1)(598)    <= not(local_tmr_voter(597));                                                                           
                tmr_registers(2)(598)    <= not(local_tmr_voter(597));                                                                           
 
                tmr_registers(0)(599)    <= not(local_tmr_voter(598));                                                                           
                tmr_registers(1)(599)    <= not(local_tmr_voter(598));                                                                           
                tmr_registers(2)(599)    <= not(local_tmr_voter(598));                                                                           
 
                tmr_registers(0)(600)    <= not(local_tmr_voter(599));                                                                           
                tmr_registers(1)(600)    <= not(local_tmr_voter(599));                                                                           
                tmr_registers(2)(600)    <= not(local_tmr_voter(599));                                                                           
 
                tmr_registers(0)(601)    <= not(local_tmr_voter(600));                                                                           
                tmr_registers(1)(601)    <= not(local_tmr_voter(600));                                                                           
                tmr_registers(2)(601)    <= not(local_tmr_voter(600));                                                                           
 
                tmr_registers(0)(602)    <= not(local_tmr_voter(601));                                                                           
                tmr_registers(1)(602)    <= not(local_tmr_voter(601));                                                                           
                tmr_registers(2)(602)    <= not(local_tmr_voter(601));                                                                           
 
                tmr_registers(0)(603)    <= not(local_tmr_voter(602));                                                                           
                tmr_registers(1)(603)    <= not(local_tmr_voter(602));                                                                           
                tmr_registers(2)(603)    <= not(local_tmr_voter(602));                                                                           
 
                tmr_registers(0)(604)    <= not(local_tmr_voter(603));                                                                           
                tmr_registers(1)(604)    <= not(local_tmr_voter(603));                                                                           
                tmr_registers(2)(604)    <= not(local_tmr_voter(603));                                                                           
 
                tmr_registers(0)(605)    <= not(local_tmr_voter(604));                                                                           
                tmr_registers(1)(605)    <= not(local_tmr_voter(604));                                                                           
                tmr_registers(2)(605)    <= not(local_tmr_voter(604));                                                                           
 
                tmr_registers(0)(606)    <= not(local_tmr_voter(605));                                                                           
                tmr_registers(1)(606)    <= not(local_tmr_voter(605));                                                                           
                tmr_registers(2)(606)    <= not(local_tmr_voter(605));                                                                           
 
                tmr_registers(0)(607)    <= not(local_tmr_voter(606));                                                                           
                tmr_registers(1)(607)    <= not(local_tmr_voter(606));                                                                           
                tmr_registers(2)(607)    <= not(local_tmr_voter(606));                                                                           
 
                tmr_registers(0)(608)    <= not(local_tmr_voter(607));                                                                           
                tmr_registers(1)(608)    <= not(local_tmr_voter(607));                                                                           
                tmr_registers(2)(608)    <= not(local_tmr_voter(607));                                                                           
 
                tmr_registers(0)(609)    <= not(local_tmr_voter(608));                                                                           
                tmr_registers(1)(609)    <= not(local_tmr_voter(608));                                                                           
                tmr_registers(2)(609)    <= not(local_tmr_voter(608));                                                                           
 
                tmr_registers(0)(610)    <= not(local_tmr_voter(609));                                                                           
                tmr_registers(1)(610)    <= not(local_tmr_voter(609));                                                                           
                tmr_registers(2)(610)    <= not(local_tmr_voter(609));                                                                           
 
                tmr_registers(0)(611)    <= not(local_tmr_voter(610));                                                                           
                tmr_registers(1)(611)    <= not(local_tmr_voter(610));                                                                           
                tmr_registers(2)(611)    <= not(local_tmr_voter(610));                                                                           
 
                tmr_registers(0)(612)    <= not(local_tmr_voter(611));                                                                           
                tmr_registers(1)(612)    <= not(local_tmr_voter(611));                                                                           
                tmr_registers(2)(612)    <= not(local_tmr_voter(611));                                                                           
 
                tmr_registers(0)(613)    <= not(local_tmr_voter(612));                                                                           
                tmr_registers(1)(613)    <= not(local_tmr_voter(612));                                                                           
                tmr_registers(2)(613)    <= not(local_tmr_voter(612));                                                                           
 
                tmr_registers(0)(614)    <= not(local_tmr_voter(613));                                                                           
                tmr_registers(1)(614)    <= not(local_tmr_voter(613));                                                                           
                tmr_registers(2)(614)    <= not(local_tmr_voter(613));                                                                           
 
                tmr_registers(0)(615)    <= not(local_tmr_voter(614));                                                                           
                tmr_registers(1)(615)    <= not(local_tmr_voter(614));                                                                           
                tmr_registers(2)(615)    <= not(local_tmr_voter(614));                                                                           
 
                tmr_registers(0)(616)    <= not(local_tmr_voter(615));                                                                           
                tmr_registers(1)(616)    <= not(local_tmr_voter(615));                                                                           
                tmr_registers(2)(616)    <= not(local_tmr_voter(615));                                                                           
 
                tmr_registers(0)(617)    <= not(local_tmr_voter(616));                                                                           
                tmr_registers(1)(617)    <= not(local_tmr_voter(616));                                                                           
                tmr_registers(2)(617)    <= not(local_tmr_voter(616));                                                                           
 
                tmr_registers(0)(618)    <= not(local_tmr_voter(617));                                                                           
                tmr_registers(1)(618)    <= not(local_tmr_voter(617));                                                                           
                tmr_registers(2)(618)    <= not(local_tmr_voter(617));                                                                           
 
                tmr_registers(0)(619)    <= not(local_tmr_voter(618));                                                                           
                tmr_registers(1)(619)    <= not(local_tmr_voter(618));                                                                           
                tmr_registers(2)(619)    <= not(local_tmr_voter(618));                                                                           
 
                tmr_registers(0)(620)    <= not(local_tmr_voter(619));                                                                           
                tmr_registers(1)(620)    <= not(local_tmr_voter(619));                                                                           
                tmr_registers(2)(620)    <= not(local_tmr_voter(619));                                                                           
 
                tmr_registers(0)(621)    <= not(local_tmr_voter(620));                                                                           
                tmr_registers(1)(621)    <= not(local_tmr_voter(620));                                                                           
                tmr_registers(2)(621)    <= not(local_tmr_voter(620));                                                                           
 
                tmr_registers(0)(622)    <= not(local_tmr_voter(621));                                                                           
                tmr_registers(1)(622)    <= not(local_tmr_voter(621));                                                                           
                tmr_registers(2)(622)    <= not(local_tmr_voter(621));                                                                           
 
                tmr_registers(0)(623)    <= not(local_tmr_voter(622));                                                                           
                tmr_registers(1)(623)    <= not(local_tmr_voter(622));                                                                           
                tmr_registers(2)(623)    <= not(local_tmr_voter(622));                                                                           
 
                tmr_registers(0)(624)    <= not(local_tmr_voter(623));                                                                           
                tmr_registers(1)(624)    <= not(local_tmr_voter(623));                                                                           
                tmr_registers(2)(624)    <= not(local_tmr_voter(623));                                                                           
 
                tmr_registers(0)(625)    <= not(local_tmr_voter(624));                                                                           
                tmr_registers(1)(625)    <= not(local_tmr_voter(624));                                                                           
                tmr_registers(2)(625)    <= not(local_tmr_voter(624));                                                                           
 
                tmr_registers(0)(626)    <= not(local_tmr_voter(625));                                                                           
                tmr_registers(1)(626)    <= not(local_tmr_voter(625));                                                                           
                tmr_registers(2)(626)    <= not(local_tmr_voter(625));                                                                           
 
                tmr_registers(0)(627)    <= not(local_tmr_voter(626));                                                                           
                tmr_registers(1)(627)    <= not(local_tmr_voter(626));                                                                           
                tmr_registers(2)(627)    <= not(local_tmr_voter(626));                                                                           
 
                tmr_registers(0)(628)    <= not(local_tmr_voter(627));                                                                           
                tmr_registers(1)(628)    <= not(local_tmr_voter(627));                                                                           
                tmr_registers(2)(628)    <= not(local_tmr_voter(627));                                                                           
 
                tmr_registers(0)(629)    <= not(local_tmr_voter(628));                                                                           
                tmr_registers(1)(629)    <= not(local_tmr_voter(628));                                                                           
                tmr_registers(2)(629)    <= not(local_tmr_voter(628));                                                                           
 
                tmr_registers(0)(630)    <= not(local_tmr_voter(629));                                                                           
                tmr_registers(1)(630)    <= not(local_tmr_voter(629));                                                                           
                tmr_registers(2)(630)    <= not(local_tmr_voter(629));                                                                           
 
                tmr_registers(0)(631)    <= not(local_tmr_voter(630));                                                                           
                tmr_registers(1)(631)    <= not(local_tmr_voter(630));                                                                           
                tmr_registers(2)(631)    <= not(local_tmr_voter(630));                                                                           
 
                tmr_registers(0)(632)    <= not(local_tmr_voter(631));                                                                           
                tmr_registers(1)(632)    <= not(local_tmr_voter(631));                                                                           
                tmr_registers(2)(632)    <= not(local_tmr_voter(631));                                                                           
 
                tmr_registers(0)(633)    <= not(local_tmr_voter(632));                                                                           
                tmr_registers(1)(633)    <= not(local_tmr_voter(632));                                                                           
                tmr_registers(2)(633)    <= not(local_tmr_voter(632));                                                                           
 
                tmr_registers(0)(634)    <= not(local_tmr_voter(633));                                                                           
                tmr_registers(1)(634)    <= not(local_tmr_voter(633));                                                                           
                tmr_registers(2)(634)    <= not(local_tmr_voter(633));                                                                           
 
                tmr_registers(0)(635)    <= not(local_tmr_voter(634));                                                                           
                tmr_registers(1)(635)    <= not(local_tmr_voter(634));                                                                           
                tmr_registers(2)(635)    <= not(local_tmr_voter(634));                                                                           
 
                tmr_registers(0)(636)    <= not(local_tmr_voter(635));                                                                           
                tmr_registers(1)(636)    <= not(local_tmr_voter(635));                                                                           
                tmr_registers(2)(636)    <= not(local_tmr_voter(635));                                                                           
 
                tmr_registers(0)(637)    <= not(local_tmr_voter(636));                                                                           
                tmr_registers(1)(637)    <= not(local_tmr_voter(636));                                                                           
                tmr_registers(2)(637)    <= not(local_tmr_voter(636));                                                                           
 
                tmr_registers(0)(638)    <= not(local_tmr_voter(637));                                                                           
                tmr_registers(1)(638)    <= not(local_tmr_voter(637));                                                                           
                tmr_registers(2)(638)    <= not(local_tmr_voter(637));                                                                           
 
                tmr_registers(0)(639)    <= not(local_tmr_voter(638));                                                                           
                tmr_registers(1)(639)    <= not(local_tmr_voter(638));                                                                           
                tmr_registers(2)(639)    <= not(local_tmr_voter(638));                                                                           
 
                tmr_registers(0)(640)    <= not(local_tmr_voter(639));                                                                           
                tmr_registers(1)(640)    <= not(local_tmr_voter(639));                                                                           
                tmr_registers(2)(640)    <= not(local_tmr_voter(639));                                                                           
 
                tmr_registers(0)(641)    <= not(local_tmr_voter(640));                                                                           
                tmr_registers(1)(641)    <= not(local_tmr_voter(640));                                                                           
                tmr_registers(2)(641)    <= not(local_tmr_voter(640));                                                                           
 
                tmr_registers(0)(642)    <= not(local_tmr_voter(641));                                                                           
                tmr_registers(1)(642)    <= not(local_tmr_voter(641));                                                                           
                tmr_registers(2)(642)    <= not(local_tmr_voter(641));                                                                           
 
                tmr_registers(0)(643)    <= not(local_tmr_voter(642));                                                                           
                tmr_registers(1)(643)    <= not(local_tmr_voter(642));                                                                           
                tmr_registers(2)(643)    <= not(local_tmr_voter(642));                                                                           
 
                tmr_registers(0)(644)    <= not(local_tmr_voter(643));                                                                           
                tmr_registers(1)(644)    <= not(local_tmr_voter(643));                                                                           
                tmr_registers(2)(644)    <= not(local_tmr_voter(643));                                                                           
 
                tmr_registers(0)(645)    <= not(local_tmr_voter(644));                                                                           
                tmr_registers(1)(645)    <= not(local_tmr_voter(644));                                                                           
                tmr_registers(2)(645)    <= not(local_tmr_voter(644));                                                                           
 
                tmr_registers(0)(646)    <= not(local_tmr_voter(645));                                                                           
                tmr_registers(1)(646)    <= not(local_tmr_voter(645));                                                                           
                tmr_registers(2)(646)    <= not(local_tmr_voter(645));                                                                           
 
                tmr_registers(0)(647)    <= not(local_tmr_voter(646));                                                                           
                tmr_registers(1)(647)    <= not(local_tmr_voter(646));                                                                           
                tmr_registers(2)(647)    <= not(local_tmr_voter(646));                                                                           
 
                tmr_registers(0)(648)    <= not(local_tmr_voter(647));                                                                           
                tmr_registers(1)(648)    <= not(local_tmr_voter(647));                                                                           
                tmr_registers(2)(648)    <= not(local_tmr_voter(647));                                                                           
 
                tmr_registers(0)(649)    <= not(local_tmr_voter(648));                                                                           
                tmr_registers(1)(649)    <= not(local_tmr_voter(648));                                                                           
                tmr_registers(2)(649)    <= not(local_tmr_voter(648));                                                                           
 
                tmr_registers(0)(650)    <= not(local_tmr_voter(649));                                                                           
                tmr_registers(1)(650)    <= not(local_tmr_voter(649));                                                                           
                tmr_registers(2)(650)    <= not(local_tmr_voter(649));                                                                           
 
                tmr_registers(0)(651)    <= not(local_tmr_voter(650));                                                                           
                tmr_registers(1)(651)    <= not(local_tmr_voter(650));                                                                           
                tmr_registers(2)(651)    <= not(local_tmr_voter(650));                                                                           
 
                tmr_registers(0)(652)    <= not(local_tmr_voter(651));                                                                           
                tmr_registers(1)(652)    <= not(local_tmr_voter(651));                                                                           
                tmr_registers(2)(652)    <= not(local_tmr_voter(651));                                                                           
 
                tmr_registers(0)(653)    <= not(local_tmr_voter(652));                                                                           
                tmr_registers(1)(653)    <= not(local_tmr_voter(652));                                                                           
                tmr_registers(2)(653)    <= not(local_tmr_voter(652));                                                                           
 
                tmr_registers(0)(654)    <= not(local_tmr_voter(653));                                                                           
                tmr_registers(1)(654)    <= not(local_tmr_voter(653));                                                                           
                tmr_registers(2)(654)    <= not(local_tmr_voter(653));                                                                           
 
                tmr_registers(0)(655)    <= not(local_tmr_voter(654));                                                                           
                tmr_registers(1)(655)    <= not(local_tmr_voter(654));                                                                           
                tmr_registers(2)(655)    <= not(local_tmr_voter(654));                                                                           
 
                tmr_registers(0)(656)    <= not(local_tmr_voter(655));                                                                           
                tmr_registers(1)(656)    <= not(local_tmr_voter(655));                                                                           
                tmr_registers(2)(656)    <= not(local_tmr_voter(655));                                                                           
 
                tmr_registers(0)(657)    <= not(local_tmr_voter(656));                                                                           
                tmr_registers(1)(657)    <= not(local_tmr_voter(656));                                                                           
                tmr_registers(2)(657)    <= not(local_tmr_voter(656));                                                                           
 
                tmr_registers(0)(658)    <= not(local_tmr_voter(657));                                                                           
                tmr_registers(1)(658)    <= not(local_tmr_voter(657));                                                                           
                tmr_registers(2)(658)    <= not(local_tmr_voter(657));                                                                           
 
                tmr_registers(0)(659)    <= not(local_tmr_voter(658));                                                                           
                tmr_registers(1)(659)    <= not(local_tmr_voter(658));                                                                           
                tmr_registers(2)(659)    <= not(local_tmr_voter(658));                                                                           
 
                tmr_registers(0)(660)    <= not(local_tmr_voter(659));                                                                           
                tmr_registers(1)(660)    <= not(local_tmr_voter(659));                                                                           
                tmr_registers(2)(660)    <= not(local_tmr_voter(659));                                                                           
 
                tmr_registers(0)(661)    <= not(local_tmr_voter(660));                                                                           
                tmr_registers(1)(661)    <= not(local_tmr_voter(660));                                                                           
                tmr_registers(2)(661)    <= not(local_tmr_voter(660));                                                                           
 
                tmr_registers(0)(662)    <= not(local_tmr_voter(661));                                                                           
                tmr_registers(1)(662)    <= not(local_tmr_voter(661));                                                                           
                tmr_registers(2)(662)    <= not(local_tmr_voter(661));                                                                           
 
                tmr_registers(0)(663)    <= not(local_tmr_voter(662));                                                                           
                tmr_registers(1)(663)    <= not(local_tmr_voter(662));                                                                           
                tmr_registers(2)(663)    <= not(local_tmr_voter(662));                                                                           
 
                tmr_registers(0)(664)    <= not(local_tmr_voter(663));                                                                           
                tmr_registers(1)(664)    <= not(local_tmr_voter(663));                                                                           
                tmr_registers(2)(664)    <= not(local_tmr_voter(663));                                                                           
 
                tmr_registers(0)(665)    <= not(local_tmr_voter(664));                                                                           
                tmr_registers(1)(665)    <= not(local_tmr_voter(664));                                                                           
                tmr_registers(2)(665)    <= not(local_tmr_voter(664));                                                                           
 
                tmr_registers(0)(666)    <= not(local_tmr_voter(665));                                                                           
                tmr_registers(1)(666)    <= not(local_tmr_voter(665));                                                                           
                tmr_registers(2)(666)    <= not(local_tmr_voter(665));                                                                           
 
                tmr_registers(0)(667)    <= not(local_tmr_voter(666));                                                                           
                tmr_registers(1)(667)    <= not(local_tmr_voter(666));                                                                           
                tmr_registers(2)(667)    <= not(local_tmr_voter(666));                                                                           
 
                tmr_registers(0)(668)    <= not(local_tmr_voter(667));                                                                           
                tmr_registers(1)(668)    <= not(local_tmr_voter(667));                                                                           
                tmr_registers(2)(668)    <= not(local_tmr_voter(667));                                                                           
 
                tmr_registers(0)(669)    <= not(local_tmr_voter(668));                                                                           
                tmr_registers(1)(669)    <= not(local_tmr_voter(668));                                                                           
                tmr_registers(2)(669)    <= not(local_tmr_voter(668));                                                                           
 
                tmr_registers(0)(670)    <= not(local_tmr_voter(669));                                                                           
                tmr_registers(1)(670)    <= not(local_tmr_voter(669));                                                                           
                tmr_registers(2)(670)    <= not(local_tmr_voter(669));                                                                           
 
                tmr_registers(0)(671)    <= not(local_tmr_voter(670));                                                                           
                tmr_registers(1)(671)    <= not(local_tmr_voter(670));                                                                           
                tmr_registers(2)(671)    <= not(local_tmr_voter(670));                                                                           
 
                tmr_registers(0)(672)    <= not(local_tmr_voter(671));                                                                           
                tmr_registers(1)(672)    <= not(local_tmr_voter(671));                                                                           
                tmr_registers(2)(672)    <= not(local_tmr_voter(671));                                                                           
 
                tmr_registers(0)(673)    <= not(local_tmr_voter(672));                                                                           
                tmr_registers(1)(673)    <= not(local_tmr_voter(672));                                                                           
                tmr_registers(2)(673)    <= not(local_tmr_voter(672));                                                                           
 
                tmr_registers(0)(674)    <= not(local_tmr_voter(673));                                                                           
                tmr_registers(1)(674)    <= not(local_tmr_voter(673));                                                                           
                tmr_registers(2)(674)    <= not(local_tmr_voter(673));                                                                           
 
                tmr_registers(0)(675)    <= not(local_tmr_voter(674));                                                                           
                tmr_registers(1)(675)    <= not(local_tmr_voter(674));                                                                           
                tmr_registers(2)(675)    <= not(local_tmr_voter(674));                                                                           
 
                tmr_registers(0)(676)    <= not(local_tmr_voter(675));                                                                           
                tmr_registers(1)(676)    <= not(local_tmr_voter(675));                                                                           
                tmr_registers(2)(676)    <= not(local_tmr_voter(675));                                                                           
 
                tmr_registers(0)(677)    <= not(local_tmr_voter(676));                                                                           
                tmr_registers(1)(677)    <= not(local_tmr_voter(676));                                                                           
                tmr_registers(2)(677)    <= not(local_tmr_voter(676));                                                                           
 
                tmr_registers(0)(678)    <= not(local_tmr_voter(677));                                                                           
                tmr_registers(1)(678)    <= not(local_tmr_voter(677));                                                                           
                tmr_registers(2)(678)    <= not(local_tmr_voter(677));                                                                           
 
                tmr_registers(0)(679)    <= not(local_tmr_voter(678));                                                                           
                tmr_registers(1)(679)    <= not(local_tmr_voter(678));                                                                           
                tmr_registers(2)(679)    <= not(local_tmr_voter(678));                                                                           
 
                tmr_registers(0)(680)    <= not(local_tmr_voter(679));                                                                           
                tmr_registers(1)(680)    <= not(local_tmr_voter(679));                                                                           
                tmr_registers(2)(680)    <= not(local_tmr_voter(679));                                                                           
 
                tmr_registers(0)(681)    <= not(local_tmr_voter(680));                                                                           
                tmr_registers(1)(681)    <= not(local_tmr_voter(680));                                                                           
                tmr_registers(2)(681)    <= not(local_tmr_voter(680));                                                                           
 
                tmr_registers(0)(682)    <= not(local_tmr_voter(681));                                                                           
                tmr_registers(1)(682)    <= not(local_tmr_voter(681));                                                                           
                tmr_registers(2)(682)    <= not(local_tmr_voter(681));                                                                           
 
                tmr_registers(0)(683)    <= not(local_tmr_voter(682));                                                                           
                tmr_registers(1)(683)    <= not(local_tmr_voter(682));                                                                           
                tmr_registers(2)(683)    <= not(local_tmr_voter(682));                                                                           
 
                tmr_registers(0)(684)    <= not(local_tmr_voter(683));                                                                           
                tmr_registers(1)(684)    <= not(local_tmr_voter(683));                                                                           
                tmr_registers(2)(684)    <= not(local_tmr_voter(683));                                                                           
 
                tmr_registers(0)(685)    <= not(local_tmr_voter(684));                                                                           
                tmr_registers(1)(685)    <= not(local_tmr_voter(684));                                                                           
                tmr_registers(2)(685)    <= not(local_tmr_voter(684));                                                                           
 
                tmr_registers(0)(686)    <= not(local_tmr_voter(685));                                                                           
                tmr_registers(1)(686)    <= not(local_tmr_voter(685));                                                                           
                tmr_registers(2)(686)    <= not(local_tmr_voter(685));                                                                           
 
                tmr_registers(0)(687)    <= not(local_tmr_voter(686));                                                                           
                tmr_registers(1)(687)    <= not(local_tmr_voter(686));                                                                           
                tmr_registers(2)(687)    <= not(local_tmr_voter(686));                                                                           
 
                tmr_registers(0)(688)    <= not(local_tmr_voter(687));                                                                           
                tmr_registers(1)(688)    <= not(local_tmr_voter(687));                                                                           
                tmr_registers(2)(688)    <= not(local_tmr_voter(687));                                                                           
 
                tmr_registers(0)(689)    <= not(local_tmr_voter(688));                                                                           
                tmr_registers(1)(689)    <= not(local_tmr_voter(688));                                                                           
                tmr_registers(2)(689)    <= not(local_tmr_voter(688));                                                                           
 
                tmr_registers(0)(690)    <= not(local_tmr_voter(689));                                                                           
                tmr_registers(1)(690)    <= not(local_tmr_voter(689));                                                                           
                tmr_registers(2)(690)    <= not(local_tmr_voter(689));                                                                           
 
                tmr_registers(0)(691)    <= not(local_tmr_voter(690));                                                                           
                tmr_registers(1)(691)    <= not(local_tmr_voter(690));                                                                           
                tmr_registers(2)(691)    <= not(local_tmr_voter(690));                                                                           
 
                tmr_registers(0)(692)    <= not(local_tmr_voter(691));                                                                           
                tmr_registers(1)(692)    <= not(local_tmr_voter(691));                                                                           
                tmr_registers(2)(692)    <= not(local_tmr_voter(691));                                                                           
 
                tmr_registers(0)(693)    <= not(local_tmr_voter(692));                                                                           
                tmr_registers(1)(693)    <= not(local_tmr_voter(692));                                                                           
                tmr_registers(2)(693)    <= not(local_tmr_voter(692));                                                                           
 
                tmr_registers(0)(694)    <= not(local_tmr_voter(693));                                                                           
                tmr_registers(1)(694)    <= not(local_tmr_voter(693));                                                                           
                tmr_registers(2)(694)    <= not(local_tmr_voter(693));                                                                           
 
                tmr_registers(0)(695)    <= not(local_tmr_voter(694));                                                                           
                tmr_registers(1)(695)    <= not(local_tmr_voter(694));                                                                           
                tmr_registers(2)(695)    <= not(local_tmr_voter(694));                                                                           
 
                tmr_registers(0)(696)    <= not(local_tmr_voter(695));                                                                           
                tmr_registers(1)(696)    <= not(local_tmr_voter(695));                                                                           
                tmr_registers(2)(696)    <= not(local_tmr_voter(695));                                                                           
 
                tmr_registers(0)(697)    <= not(local_tmr_voter(696));                                                                           
                tmr_registers(1)(697)    <= not(local_tmr_voter(696));                                                                           
                tmr_registers(2)(697)    <= not(local_tmr_voter(696));                                                                           
 
                tmr_registers(0)(698)    <= not(local_tmr_voter(697));                                                                           
                tmr_registers(1)(698)    <= not(local_tmr_voter(697));                                                                           
                tmr_registers(2)(698)    <= not(local_tmr_voter(697));                                                                           
 
                tmr_registers(0)(699)    <= not(local_tmr_voter(698));                                                                           
                tmr_registers(1)(699)    <= not(local_tmr_voter(698));                                                                           
                tmr_registers(2)(699)    <= not(local_tmr_voter(698));                                                                           
 
                tmr_registers(0)(700)    <= not(local_tmr_voter(699));                                                                           
                tmr_registers(1)(700)    <= not(local_tmr_voter(699));                                                                           
                tmr_registers(2)(700)    <= not(local_tmr_voter(699));                                                                           
 
                tmr_registers(0)(701)    <= not(local_tmr_voter(700));                                                                           
                tmr_registers(1)(701)    <= not(local_tmr_voter(700));                                                                           
                tmr_registers(2)(701)    <= not(local_tmr_voter(700));                                                                           
 
                tmr_registers(0)(702)    <= not(local_tmr_voter(701));                                                                           
                tmr_registers(1)(702)    <= not(local_tmr_voter(701));                                                                           
                tmr_registers(2)(702)    <= not(local_tmr_voter(701));                                                                           
 
                tmr_registers(0)(703)    <= not(local_tmr_voter(702));                                                                           
                tmr_registers(1)(703)    <= not(local_tmr_voter(702));                                                                           
                tmr_registers(2)(703)    <= not(local_tmr_voter(702));                                                                           
 
                tmr_registers(0)(704)    <= not(local_tmr_voter(703));                                                                           
                tmr_registers(1)(704)    <= not(local_tmr_voter(703));                                                                           
                tmr_registers(2)(704)    <= not(local_tmr_voter(703));                                                                           
 
                tmr_registers(0)(705)    <= not(local_tmr_voter(704));                                                                           
                tmr_registers(1)(705)    <= not(local_tmr_voter(704));                                                                           
                tmr_registers(2)(705)    <= not(local_tmr_voter(704));                                                                           
 
                tmr_registers(0)(706)    <= not(local_tmr_voter(705));                                                                           
                tmr_registers(1)(706)    <= not(local_tmr_voter(705));                                                                           
                tmr_registers(2)(706)    <= not(local_tmr_voter(705));                                                                           
 
                tmr_registers(0)(707)    <= not(local_tmr_voter(706));                                                                           
                tmr_registers(1)(707)    <= not(local_tmr_voter(706));                                                                           
                tmr_registers(2)(707)    <= not(local_tmr_voter(706));                                                                           
 
                tmr_registers(0)(708)    <= not(local_tmr_voter(707));                                                                           
                tmr_registers(1)(708)    <= not(local_tmr_voter(707));                                                                           
                tmr_registers(2)(708)    <= not(local_tmr_voter(707));                                                                           
 
                tmr_registers(0)(709)    <= not(local_tmr_voter(708));                                                                           
                tmr_registers(1)(709)    <= not(local_tmr_voter(708));                                                                           
                tmr_registers(2)(709)    <= not(local_tmr_voter(708));                                                                           
 
                tmr_registers(0)(710)    <= not(local_tmr_voter(709));                                                                           
                tmr_registers(1)(710)    <= not(local_tmr_voter(709));                                                                           
                tmr_registers(2)(710)    <= not(local_tmr_voter(709));                                                                           
 
                tmr_registers(0)(711)    <= not(local_tmr_voter(710));                                                                           
                tmr_registers(1)(711)    <= not(local_tmr_voter(710));                                                                           
                tmr_registers(2)(711)    <= not(local_tmr_voter(710));                                                                           
 
                tmr_registers(0)(712)    <= not(local_tmr_voter(711));                                                                           
                tmr_registers(1)(712)    <= not(local_tmr_voter(711));                                                                           
                tmr_registers(2)(712)    <= not(local_tmr_voter(711));                                                                           
 
                tmr_registers(0)(713)    <= not(local_tmr_voter(712));                                                                           
                tmr_registers(1)(713)    <= not(local_tmr_voter(712));                                                                           
                tmr_registers(2)(713)    <= not(local_tmr_voter(712));                                                                           
 
                tmr_registers(0)(714)    <= not(local_tmr_voter(713));                                                                           
                tmr_registers(1)(714)    <= not(local_tmr_voter(713));                                                                           
                tmr_registers(2)(714)    <= not(local_tmr_voter(713));                                                                           
 
                tmr_registers(0)(715)    <= not(local_tmr_voter(714));                                                                           
                tmr_registers(1)(715)    <= not(local_tmr_voter(714));                                                                           
                tmr_registers(2)(715)    <= not(local_tmr_voter(714));                                                                           
 
                tmr_registers(0)(716)    <= not(local_tmr_voter(715));                                                                           
                tmr_registers(1)(716)    <= not(local_tmr_voter(715));                                                                           
                tmr_registers(2)(716)    <= not(local_tmr_voter(715));                                                                           
 
                tmr_registers(0)(717)    <= not(local_tmr_voter(716));                                                                           
                tmr_registers(1)(717)    <= not(local_tmr_voter(716));                                                                           
                tmr_registers(2)(717)    <= not(local_tmr_voter(716));                                                                           
 
                tmr_registers(0)(718)    <= not(local_tmr_voter(717));                                                                           
                tmr_registers(1)(718)    <= not(local_tmr_voter(717));                                                                           
                tmr_registers(2)(718)    <= not(local_tmr_voter(717));                                                                           
 
                tmr_registers(0)(719)    <= not(local_tmr_voter(718));                                                                           
                tmr_registers(1)(719)    <= not(local_tmr_voter(718));                                                                           
                tmr_registers(2)(719)    <= not(local_tmr_voter(718));                                                                           
 
                tmr_registers(0)(720)    <= not(local_tmr_voter(719));                                                                           
                tmr_registers(1)(720)    <= not(local_tmr_voter(719));                                                                           
                tmr_registers(2)(720)    <= not(local_tmr_voter(719));                                                                           
 
                tmr_registers(0)(721)    <= not(local_tmr_voter(720));                                                                           
                tmr_registers(1)(721)    <= not(local_tmr_voter(720));                                                                           
                tmr_registers(2)(721)    <= not(local_tmr_voter(720));                                                                           
 
                tmr_registers(0)(722)    <= not(local_tmr_voter(721));                                                                           
                tmr_registers(1)(722)    <= not(local_tmr_voter(721));                                                                           
                tmr_registers(2)(722)    <= not(local_tmr_voter(721));                                                                           
 
                tmr_registers(0)(723)    <= not(local_tmr_voter(722));                                                                           
                tmr_registers(1)(723)    <= not(local_tmr_voter(722));                                                                           
                tmr_registers(2)(723)    <= not(local_tmr_voter(722));                                                                           
 
                tmr_registers(0)(724)    <= not(local_tmr_voter(723));                                                                           
                tmr_registers(1)(724)    <= not(local_tmr_voter(723));                                                                           
                tmr_registers(2)(724)    <= not(local_tmr_voter(723));                                                                           
 
                tmr_registers(0)(725)    <= not(local_tmr_voter(724));                                                                           
                tmr_registers(1)(725)    <= not(local_tmr_voter(724));                                                                           
                tmr_registers(2)(725)    <= not(local_tmr_voter(724));                                                                           
 
                tmr_registers(0)(726)    <= not(local_tmr_voter(725));                                                                           
                tmr_registers(1)(726)    <= not(local_tmr_voter(725));                                                                           
                tmr_registers(2)(726)    <= not(local_tmr_voter(725));                                                                           
 
                tmr_registers(0)(727)    <= not(local_tmr_voter(726));                                                                           
                tmr_registers(1)(727)    <= not(local_tmr_voter(726));                                                                           
                tmr_registers(2)(727)    <= not(local_tmr_voter(726));                                                                           
 
                tmr_registers(0)(728)    <= not(local_tmr_voter(727));                                                                           
                tmr_registers(1)(728)    <= not(local_tmr_voter(727));                                                                           
                tmr_registers(2)(728)    <= not(local_tmr_voter(727));                                                                           
 
                tmr_registers(0)(729)    <= not(local_tmr_voter(728));                                                                           
                tmr_registers(1)(729)    <= not(local_tmr_voter(728));                                                                           
                tmr_registers(2)(729)    <= not(local_tmr_voter(728));                                                                           
 
                tmr_registers(0)(730)    <= not(local_tmr_voter(729));                                                                           
                tmr_registers(1)(730)    <= not(local_tmr_voter(729));                                                                           
                tmr_registers(2)(730)    <= not(local_tmr_voter(729));                                                                           
 
                tmr_registers(0)(731)    <= not(local_tmr_voter(730));                                                                           
                tmr_registers(1)(731)    <= not(local_tmr_voter(730));                                                                           
                tmr_registers(2)(731)    <= not(local_tmr_voter(730));                                                                           
 
                tmr_registers(0)(732)    <= not(local_tmr_voter(731));                                                                           
                tmr_registers(1)(732)    <= not(local_tmr_voter(731));                                                                           
                tmr_registers(2)(732)    <= not(local_tmr_voter(731));                                                                           
 
                tmr_registers(0)(733)    <= not(local_tmr_voter(732));                                                                           
                tmr_registers(1)(733)    <= not(local_tmr_voter(732));                                                                           
                tmr_registers(2)(733)    <= not(local_tmr_voter(732));                                                                           
 
                tmr_registers(0)(734)    <= not(local_tmr_voter(733));                                                                           
                tmr_registers(1)(734)    <= not(local_tmr_voter(733));                                                                           
                tmr_registers(2)(734)    <= not(local_tmr_voter(733));                                                                           
 
                tmr_registers(0)(735)    <= not(local_tmr_voter(734));                                                                           
                tmr_registers(1)(735)    <= not(local_tmr_voter(734));                                                                           
                tmr_registers(2)(735)    <= not(local_tmr_voter(734));                                                                           
 
                tmr_registers(0)(736)    <= not(local_tmr_voter(735));                                                                           
                tmr_registers(1)(736)    <= not(local_tmr_voter(735));                                                                           
                tmr_registers(2)(736)    <= not(local_tmr_voter(735));                                                                           
 
                tmr_registers(0)(737)    <= not(local_tmr_voter(736));                                                                           
                tmr_registers(1)(737)    <= not(local_tmr_voter(736));                                                                           
                tmr_registers(2)(737)    <= not(local_tmr_voter(736));                                                                           
 
                tmr_registers(0)(738)    <= not(local_tmr_voter(737));                                                                           
                tmr_registers(1)(738)    <= not(local_tmr_voter(737));                                                                           
                tmr_registers(2)(738)    <= not(local_tmr_voter(737));                                                                           
 
                tmr_registers(0)(739)    <= not(local_tmr_voter(738));                                                                           
                tmr_registers(1)(739)    <= not(local_tmr_voter(738));                                                                           
                tmr_registers(2)(739)    <= not(local_tmr_voter(738));                                                                           
 
                tmr_registers(0)(740)    <= not(local_tmr_voter(739));                                                                           
                tmr_registers(1)(740)    <= not(local_tmr_voter(739));                                                                           
                tmr_registers(2)(740)    <= not(local_tmr_voter(739));                                                                           
 
                tmr_registers(0)(741)    <= not(local_tmr_voter(740));                                                                           
                tmr_registers(1)(741)    <= not(local_tmr_voter(740));                                                                           
                tmr_registers(2)(741)    <= not(local_tmr_voter(740));                                                                           
 
                tmr_registers(0)(742)    <= not(local_tmr_voter(741));                                                                           
                tmr_registers(1)(742)    <= not(local_tmr_voter(741));                                                                           
                tmr_registers(2)(742)    <= not(local_tmr_voter(741));                                                                           
 
                tmr_registers(0)(743)    <= not(local_tmr_voter(742));                                                                           
                tmr_registers(1)(743)    <= not(local_tmr_voter(742));                                                                           
                tmr_registers(2)(743)    <= not(local_tmr_voter(742));                                                                           
 
                tmr_registers(0)(744)    <= not(local_tmr_voter(743));                                                                           
                tmr_registers(1)(744)    <= not(local_tmr_voter(743));                                                                           
                tmr_registers(2)(744)    <= not(local_tmr_voter(743));                                                                           
 
                tmr_registers(0)(745)    <= not(local_tmr_voter(744));                                                                           
                tmr_registers(1)(745)    <= not(local_tmr_voter(744));                                                                           
                tmr_registers(2)(745)    <= not(local_tmr_voter(744));                                                                           
 
                tmr_registers(0)(746)    <= not(local_tmr_voter(745));                                                                           
                tmr_registers(1)(746)    <= not(local_tmr_voter(745));                                                                           
                tmr_registers(2)(746)    <= not(local_tmr_voter(745));                                                                           
 
                tmr_registers(0)(747)    <= not(local_tmr_voter(746));                                                                           
                tmr_registers(1)(747)    <= not(local_tmr_voter(746));                                                                           
                tmr_registers(2)(747)    <= not(local_tmr_voter(746));                                                                           
 
                tmr_registers(0)(748)    <= not(local_tmr_voter(747));                                                                           
                tmr_registers(1)(748)    <= not(local_tmr_voter(747));                                                                           
                tmr_registers(2)(748)    <= not(local_tmr_voter(747));                                                                           
 
                tmr_registers(0)(749)    <= not(local_tmr_voter(748));                                                                           
                tmr_registers(1)(749)    <= not(local_tmr_voter(748));                                                                           
                tmr_registers(2)(749)    <= not(local_tmr_voter(748));                                                                           
 
                tmr_registers(0)(750)    <= not(local_tmr_voter(749));                                                                           
                tmr_registers(1)(750)    <= not(local_tmr_voter(749));                                                                           
                tmr_registers(2)(750)    <= not(local_tmr_voter(749));                                                                           
 
                tmr_registers(0)(751)    <= not(local_tmr_voter(750));                                                                           
                tmr_registers(1)(751)    <= not(local_tmr_voter(750));                                                                           
                tmr_registers(2)(751)    <= not(local_tmr_voter(750));                                                                           
 
                tmr_registers(0)(752)    <= not(local_tmr_voter(751));                                                                           
                tmr_registers(1)(752)    <= not(local_tmr_voter(751));                                                                           
                tmr_registers(2)(752)    <= not(local_tmr_voter(751));                                                                           
 
                tmr_registers(0)(753)    <= not(local_tmr_voter(752));                                                                           
                tmr_registers(1)(753)    <= not(local_tmr_voter(752));                                                                           
                tmr_registers(2)(753)    <= not(local_tmr_voter(752));                                                                           
 
                tmr_registers(0)(754)    <= not(local_tmr_voter(753));                                                                           
                tmr_registers(1)(754)    <= not(local_tmr_voter(753));                                                                           
                tmr_registers(2)(754)    <= not(local_tmr_voter(753));                                                                           
 
                tmr_registers(0)(755)    <= not(local_tmr_voter(754));                                                                           
                tmr_registers(1)(755)    <= not(local_tmr_voter(754));                                                                           
                tmr_registers(2)(755)    <= not(local_tmr_voter(754));                                                                           
 
                tmr_registers(0)(756)    <= not(local_tmr_voter(755));                                                                           
                tmr_registers(1)(756)    <= not(local_tmr_voter(755));                                                                           
                tmr_registers(2)(756)    <= not(local_tmr_voter(755));                                                                           
 
                tmr_registers(0)(757)    <= not(local_tmr_voter(756));                                                                           
                tmr_registers(1)(757)    <= not(local_tmr_voter(756));                                                                           
                tmr_registers(2)(757)    <= not(local_tmr_voter(756));                                                                           
 
                tmr_registers(0)(758)    <= not(local_tmr_voter(757));                                                                           
                tmr_registers(1)(758)    <= not(local_tmr_voter(757));                                                                           
                tmr_registers(2)(758)    <= not(local_tmr_voter(757));                                                                           
 
                tmr_registers(0)(759)    <= not(local_tmr_voter(758));                                                                           
                tmr_registers(1)(759)    <= not(local_tmr_voter(758));                                                                           
                tmr_registers(2)(759)    <= not(local_tmr_voter(758));                                                                           
 
                tmr_registers(0)(760)    <= not(local_tmr_voter(759));                                                                           
                tmr_registers(1)(760)    <= not(local_tmr_voter(759));                                                                           
                tmr_registers(2)(760)    <= not(local_tmr_voter(759));                                                                           
 
                tmr_registers(0)(761)    <= not(local_tmr_voter(760));                                                                           
                tmr_registers(1)(761)    <= not(local_tmr_voter(760));                                                                           
                tmr_registers(2)(761)    <= not(local_tmr_voter(760));                                                                           
 
                tmr_registers(0)(762)    <= not(local_tmr_voter(761));                                                                           
                tmr_registers(1)(762)    <= not(local_tmr_voter(761));                                                                           
                tmr_registers(2)(762)    <= not(local_tmr_voter(761));                                                                           
 
                tmr_registers(0)(763)    <= not(local_tmr_voter(762));                                                                           
                tmr_registers(1)(763)    <= not(local_tmr_voter(762));                                                                           
                tmr_registers(2)(763)    <= not(local_tmr_voter(762));                                                                           
 
                tmr_registers(0)(764)    <= not(local_tmr_voter(763));                                                                           
                tmr_registers(1)(764)    <= not(local_tmr_voter(763));                                                                           
                tmr_registers(2)(764)    <= not(local_tmr_voter(763));                                                                           
 
                tmr_registers(0)(765)    <= not(local_tmr_voter(764));                                                                           
                tmr_registers(1)(765)    <= not(local_tmr_voter(764));                                                                           
                tmr_registers(2)(765)    <= not(local_tmr_voter(764));                                                                           
 
                tmr_registers(0)(766)    <= not(local_tmr_voter(765));                                                                           
                tmr_registers(1)(766)    <= not(local_tmr_voter(765));                                                                           
                tmr_registers(2)(766)    <= not(local_tmr_voter(765));                                                                           
 
                tmr_registers(0)(767)    <= not(local_tmr_voter(766));                                                                           
                tmr_registers(1)(767)    <= not(local_tmr_voter(766));                                                                           
                tmr_registers(2)(767)    <= not(local_tmr_voter(766));                                                                           
 
                tmr_registers(0)(768)    <= not(local_tmr_voter(767));                                                                           
                tmr_registers(1)(768)    <= not(local_tmr_voter(767));                                                                           
                tmr_registers(2)(768)    <= not(local_tmr_voter(767));                                                                           
 
                tmr_registers(0)(769)    <= not(local_tmr_voter(768));                                                                           
                tmr_registers(1)(769)    <= not(local_tmr_voter(768));                                                                           
                tmr_registers(2)(769)    <= not(local_tmr_voter(768));                                                                           
 
                tmr_registers(0)(770)    <= not(local_tmr_voter(769));                                                                           
                tmr_registers(1)(770)    <= not(local_tmr_voter(769));                                                                           
                tmr_registers(2)(770)    <= not(local_tmr_voter(769));                                                                           
 
                tmr_registers(0)(771)    <= not(local_tmr_voter(770));                                                                           
                tmr_registers(1)(771)    <= not(local_tmr_voter(770));                                                                           
                tmr_registers(2)(771)    <= not(local_tmr_voter(770));                                                                           
 
                tmr_registers(0)(772)    <= not(local_tmr_voter(771));                                                                           
                tmr_registers(1)(772)    <= not(local_tmr_voter(771));                                                                           
                tmr_registers(2)(772)    <= not(local_tmr_voter(771));                                                                           
 
                tmr_registers(0)(773)    <= not(local_tmr_voter(772));                                                                           
                tmr_registers(1)(773)    <= not(local_tmr_voter(772));                                                                           
                tmr_registers(2)(773)    <= not(local_tmr_voter(772));                                                                           
 
                tmr_registers(0)(774)    <= not(local_tmr_voter(773));                                                                           
                tmr_registers(1)(774)    <= not(local_tmr_voter(773));                                                                           
                tmr_registers(2)(774)    <= not(local_tmr_voter(773));                                                                           
 
                tmr_registers(0)(775)    <= not(local_tmr_voter(774));                                                                           
                tmr_registers(1)(775)    <= not(local_tmr_voter(774));                                                                           
                tmr_registers(2)(775)    <= not(local_tmr_voter(774));                                                                           
 
                tmr_registers(0)(776)    <= not(local_tmr_voter(775));                                                                           
                tmr_registers(1)(776)    <= not(local_tmr_voter(775));                                                                           
                tmr_registers(2)(776)    <= not(local_tmr_voter(775));                                                                           
 
                tmr_registers(0)(777)    <= not(local_tmr_voter(776));                                                                           
                tmr_registers(1)(777)    <= not(local_tmr_voter(776));                                                                           
                tmr_registers(2)(777)    <= not(local_tmr_voter(776));                                                                           
 
                tmr_registers(0)(778)    <= not(local_tmr_voter(777));                                                                           
                tmr_registers(1)(778)    <= not(local_tmr_voter(777));                                                                           
                tmr_registers(2)(778)    <= not(local_tmr_voter(777));                                                                           
 
                tmr_registers(0)(779)    <= not(local_tmr_voter(778));                                                                           
                tmr_registers(1)(779)    <= not(local_tmr_voter(778));                                                                           
                tmr_registers(2)(779)    <= not(local_tmr_voter(778));                                                                           
 
                tmr_registers(0)(780)    <= not(local_tmr_voter(779));                                                                           
                tmr_registers(1)(780)    <= not(local_tmr_voter(779));                                                                           
                tmr_registers(2)(780)    <= not(local_tmr_voter(779));                                                                           
 
                tmr_registers(0)(781)    <= not(local_tmr_voter(780));                                                                           
                tmr_registers(1)(781)    <= not(local_tmr_voter(780));                                                                           
                tmr_registers(2)(781)    <= not(local_tmr_voter(780));                                                                           
 
                tmr_registers(0)(782)    <= not(local_tmr_voter(781));                                                                           
                tmr_registers(1)(782)    <= not(local_tmr_voter(781));                                                                           
                tmr_registers(2)(782)    <= not(local_tmr_voter(781));                                                                           
 
                tmr_registers(0)(783)    <= not(local_tmr_voter(782));                                                                           
                tmr_registers(1)(783)    <= not(local_tmr_voter(782));                                                                           
                tmr_registers(2)(783)    <= not(local_tmr_voter(782));                                                                           
 
                tmr_registers(0)(784)    <= not(local_tmr_voter(783));                                                                           
                tmr_registers(1)(784)    <= not(local_tmr_voter(783));                                                                           
                tmr_registers(2)(784)    <= not(local_tmr_voter(783));                                                                           
 
                tmr_registers(0)(785)    <= not(local_tmr_voter(784));                                                                           
                tmr_registers(1)(785)    <= not(local_tmr_voter(784));                                                                           
                tmr_registers(2)(785)    <= not(local_tmr_voter(784));                                                                           
 
                tmr_registers(0)(786)    <= not(local_tmr_voter(785));                                                                           
                tmr_registers(1)(786)    <= not(local_tmr_voter(785));                                                                           
                tmr_registers(2)(786)    <= not(local_tmr_voter(785));                                                                           
 
                tmr_registers(0)(787)    <= not(local_tmr_voter(786));                                                                           
                tmr_registers(1)(787)    <= not(local_tmr_voter(786));                                                                           
                tmr_registers(2)(787)    <= not(local_tmr_voter(786));                                                                           
 
                tmr_registers(0)(788)    <= not(local_tmr_voter(787));                                                                           
                tmr_registers(1)(788)    <= not(local_tmr_voter(787));                                                                           
                tmr_registers(2)(788)    <= not(local_tmr_voter(787));                                                                           
 
                tmr_registers(0)(789)    <= not(local_tmr_voter(788));                                                                           
                tmr_registers(1)(789)    <= not(local_tmr_voter(788));                                                                           
                tmr_registers(2)(789)    <= not(local_tmr_voter(788));                                                                           
 
                tmr_registers(0)(790)    <= not(local_tmr_voter(789));                                                                           
                tmr_registers(1)(790)    <= not(local_tmr_voter(789));                                                                           
                tmr_registers(2)(790)    <= not(local_tmr_voter(789));                                                                           
 
                tmr_registers(0)(791)    <= not(local_tmr_voter(790));                                                                           
                tmr_registers(1)(791)    <= not(local_tmr_voter(790));                                                                           
                tmr_registers(2)(791)    <= not(local_tmr_voter(790));                                                                           
 
                tmr_registers(0)(792)    <= not(local_tmr_voter(791));                                                                           
                tmr_registers(1)(792)    <= not(local_tmr_voter(791));                                                                           
                tmr_registers(2)(792)    <= not(local_tmr_voter(791));                                                                           
 
                tmr_registers(0)(793)    <= not(local_tmr_voter(792));                                                                           
                tmr_registers(1)(793)    <= not(local_tmr_voter(792));                                                                           
                tmr_registers(2)(793)    <= not(local_tmr_voter(792));                                                                           
 
                tmr_registers(0)(794)    <= not(local_tmr_voter(793));                                                                           
                tmr_registers(1)(794)    <= not(local_tmr_voter(793));                                                                           
                tmr_registers(2)(794)    <= not(local_tmr_voter(793));                                                                           
 
                tmr_registers(0)(795)    <= not(local_tmr_voter(794));                                                                           
                tmr_registers(1)(795)    <= not(local_tmr_voter(794));                                                                           
                tmr_registers(2)(795)    <= not(local_tmr_voter(794));                                                                           
 
                tmr_registers(0)(796)    <= not(local_tmr_voter(795));                                                                           
                tmr_registers(1)(796)    <= not(local_tmr_voter(795));                                                                           
                tmr_registers(2)(796)    <= not(local_tmr_voter(795));                                                                           
 
                tmr_registers(0)(797)    <= not(local_tmr_voter(796));                                                                           
                tmr_registers(1)(797)    <= not(local_tmr_voter(796));                                                                           
                tmr_registers(2)(797)    <= not(local_tmr_voter(796));                                                                           
 
                tmr_registers(0)(798)    <= not(local_tmr_voter(797));                                                                           
                tmr_registers(1)(798)    <= not(local_tmr_voter(797));                                                                           
                tmr_registers(2)(798)    <= not(local_tmr_voter(797));                                                                           
 
                tmr_registers(0)(799)    <= not(local_tmr_voter(798));                                                                           
                tmr_registers(1)(799)    <= not(local_tmr_voter(798));                                                                           
                tmr_registers(2)(799)    <= not(local_tmr_voter(798));                                                                           
 
                tmr_registers(0)(800)    <= not(local_tmr_voter(799));                                                                           
                tmr_registers(1)(800)    <= not(local_tmr_voter(799));                                                                           
                tmr_registers(2)(800)    <= not(local_tmr_voter(799));                                                                           
 
                tmr_registers(0)(801)    <= not(local_tmr_voter(800));                                                                           
                tmr_registers(1)(801)    <= not(local_tmr_voter(800));                                                                           
                tmr_registers(2)(801)    <= not(local_tmr_voter(800));                                                                           
 
                tmr_registers(0)(802)    <= not(local_tmr_voter(801));                                                                           
                tmr_registers(1)(802)    <= not(local_tmr_voter(801));                                                                           
                tmr_registers(2)(802)    <= not(local_tmr_voter(801));                                                                           
 
                tmr_registers(0)(803)    <= not(local_tmr_voter(802));                                                                           
                tmr_registers(1)(803)    <= not(local_tmr_voter(802));                                                                           
                tmr_registers(2)(803)    <= not(local_tmr_voter(802));                                                                           
 
                tmr_registers(0)(804)    <= not(local_tmr_voter(803));                                                                           
                tmr_registers(1)(804)    <= not(local_tmr_voter(803));                                                                           
                tmr_registers(2)(804)    <= not(local_tmr_voter(803));                                                                           
 
                tmr_registers(0)(805)    <= not(local_tmr_voter(804));                                                                           
                tmr_registers(1)(805)    <= not(local_tmr_voter(804));                                                                           
                tmr_registers(2)(805)    <= not(local_tmr_voter(804));                                                                           
 
                tmr_registers(0)(806)    <= not(local_tmr_voter(805));                                                                           
                tmr_registers(1)(806)    <= not(local_tmr_voter(805));                                                                           
                tmr_registers(2)(806)    <= not(local_tmr_voter(805));                                                                           
 
                tmr_registers(0)(807)    <= not(local_tmr_voter(806));                                                                           
                tmr_registers(1)(807)    <= not(local_tmr_voter(806));                                                                           
                tmr_registers(2)(807)    <= not(local_tmr_voter(806));                                                                           
 
                tmr_registers(0)(808)    <= not(local_tmr_voter(807));                                                                           
                tmr_registers(1)(808)    <= not(local_tmr_voter(807));                                                                           
                tmr_registers(2)(808)    <= not(local_tmr_voter(807));                                                                           
 
                tmr_registers(0)(809)    <= not(local_tmr_voter(808));                                                                           
                tmr_registers(1)(809)    <= not(local_tmr_voter(808));                                                                           
                tmr_registers(2)(809)    <= not(local_tmr_voter(808));                                                                           
 
                tmr_registers(0)(810)    <= not(local_tmr_voter(809));                                                                           
                tmr_registers(1)(810)    <= not(local_tmr_voter(809));                                                                           
                tmr_registers(2)(810)    <= not(local_tmr_voter(809));                                                                           
 
                tmr_registers(0)(811)    <= not(local_tmr_voter(810));                                                                           
                tmr_registers(1)(811)    <= not(local_tmr_voter(810));                                                                           
                tmr_registers(2)(811)    <= not(local_tmr_voter(810));                                                                           
 
                tmr_registers(0)(812)    <= not(local_tmr_voter(811));                                                                           
                tmr_registers(1)(812)    <= not(local_tmr_voter(811));                                                                           
                tmr_registers(2)(812)    <= not(local_tmr_voter(811));                                                                           
 
                tmr_registers(0)(813)    <= not(local_tmr_voter(812));                                                                           
                tmr_registers(1)(813)    <= not(local_tmr_voter(812));                                                                           
                tmr_registers(2)(813)    <= not(local_tmr_voter(812));                                                                           
 
                tmr_registers(0)(814)    <= not(local_tmr_voter(813));                                                                           
                tmr_registers(1)(814)    <= not(local_tmr_voter(813));                                                                           
                tmr_registers(2)(814)    <= not(local_tmr_voter(813));                                                                           
 
                tmr_registers(0)(815)    <= not(local_tmr_voter(814));                                                                           
                tmr_registers(1)(815)    <= not(local_tmr_voter(814));                                                                           
                tmr_registers(2)(815)    <= not(local_tmr_voter(814));                                                                           
 
                tmr_registers(0)(816)    <= not(local_tmr_voter(815));                                                                           
                tmr_registers(1)(816)    <= not(local_tmr_voter(815));                                                                           
                tmr_registers(2)(816)    <= not(local_tmr_voter(815));                                                                           
 
                tmr_registers(0)(817)    <= not(local_tmr_voter(816));                                                                           
                tmr_registers(1)(817)    <= not(local_tmr_voter(816));                                                                           
                tmr_registers(2)(817)    <= not(local_tmr_voter(816));                                                                           
 
                tmr_registers(0)(818)    <= not(local_tmr_voter(817));                                                                           
                tmr_registers(1)(818)    <= not(local_tmr_voter(817));                                                                           
                tmr_registers(2)(818)    <= not(local_tmr_voter(817));                                                                           
 
                tmr_registers(0)(819)    <= not(local_tmr_voter(818));                                                                           
                tmr_registers(1)(819)    <= not(local_tmr_voter(818));                                                                           
                tmr_registers(2)(819)    <= not(local_tmr_voter(818));                                                                           
 
                tmr_registers(0)(820)    <= not(local_tmr_voter(819));                                                                           
                tmr_registers(1)(820)    <= not(local_tmr_voter(819));                                                                           
                tmr_registers(2)(820)    <= not(local_tmr_voter(819));                                                                           
 
                tmr_registers(0)(821)    <= not(local_tmr_voter(820));                                                                           
                tmr_registers(1)(821)    <= not(local_tmr_voter(820));                                                                           
                tmr_registers(2)(821)    <= not(local_tmr_voter(820));                                                                           
 
                tmr_registers(0)(822)    <= not(local_tmr_voter(821));                                                                           
                tmr_registers(1)(822)    <= not(local_tmr_voter(821));                                                                           
                tmr_registers(2)(822)    <= not(local_tmr_voter(821));                                                                           
 
                tmr_registers(0)(823)    <= not(local_tmr_voter(822));                                                                           
                tmr_registers(1)(823)    <= not(local_tmr_voter(822));                                                                           
                tmr_registers(2)(823)    <= not(local_tmr_voter(822));                                                                           
 
                tmr_registers(0)(824)    <= not(local_tmr_voter(823));                                                                           
                tmr_registers(1)(824)    <= not(local_tmr_voter(823));                                                                           
                tmr_registers(2)(824)    <= not(local_tmr_voter(823));                                                                           
 
                tmr_registers(0)(825)    <= not(local_tmr_voter(824));                                                                           
                tmr_registers(1)(825)    <= not(local_tmr_voter(824));                                                                           
                tmr_registers(2)(825)    <= not(local_tmr_voter(824));                                                                           
 
                tmr_registers(0)(826)    <= not(local_tmr_voter(825));                                                                           
                tmr_registers(1)(826)    <= not(local_tmr_voter(825));                                                                           
                tmr_registers(2)(826)    <= not(local_tmr_voter(825));                                                                           
 
                tmr_registers(0)(827)    <= not(local_tmr_voter(826));                                                                           
                tmr_registers(1)(827)    <= not(local_tmr_voter(826));                                                                           
                tmr_registers(2)(827)    <= not(local_tmr_voter(826));                                                                           
 
                tmr_registers(0)(828)    <= not(local_tmr_voter(827));                                                                           
                tmr_registers(1)(828)    <= not(local_tmr_voter(827));                                                                           
                tmr_registers(2)(828)    <= not(local_tmr_voter(827));                                                                           
 
                tmr_registers(0)(829)    <= not(local_tmr_voter(828));                                                                           
                tmr_registers(1)(829)    <= not(local_tmr_voter(828));                                                                           
                tmr_registers(2)(829)    <= not(local_tmr_voter(828));                                                                           
 
                tmr_registers(0)(830)    <= not(local_tmr_voter(829));                                                                           
                tmr_registers(1)(830)    <= not(local_tmr_voter(829));                                                                           
                tmr_registers(2)(830)    <= not(local_tmr_voter(829));                                                                           
 
                tmr_registers(0)(831)    <= not(local_tmr_voter(830));                                                                           
                tmr_registers(1)(831)    <= not(local_tmr_voter(830));                                                                           
                tmr_registers(2)(831)    <= not(local_tmr_voter(830));                                                                           
 
                tmr_registers(0)(832)    <= not(local_tmr_voter(831));                                                                           
                tmr_registers(1)(832)    <= not(local_tmr_voter(831));                                                                           
                tmr_registers(2)(832)    <= not(local_tmr_voter(831));                                                                           
 
                tmr_registers(0)(833)    <= not(local_tmr_voter(832));                                                                           
                tmr_registers(1)(833)    <= not(local_tmr_voter(832));                                                                           
                tmr_registers(2)(833)    <= not(local_tmr_voter(832));                                                                           
 
                tmr_registers(0)(834)    <= not(local_tmr_voter(833));                                                                           
                tmr_registers(1)(834)    <= not(local_tmr_voter(833));                                                                           
                tmr_registers(2)(834)    <= not(local_tmr_voter(833));                                                                           
 
                tmr_registers(0)(835)    <= not(local_tmr_voter(834));                                                                           
                tmr_registers(1)(835)    <= not(local_tmr_voter(834));                                                                           
                tmr_registers(2)(835)    <= not(local_tmr_voter(834));                                                                           
 
                tmr_registers(0)(836)    <= not(local_tmr_voter(835));                                                                           
                tmr_registers(1)(836)    <= not(local_tmr_voter(835));                                                                           
                tmr_registers(2)(836)    <= not(local_tmr_voter(835));                                                                           
 
                tmr_registers(0)(837)    <= not(local_tmr_voter(836));                                                                           
                tmr_registers(1)(837)    <= not(local_tmr_voter(836));                                                                           
                tmr_registers(2)(837)    <= not(local_tmr_voter(836));                                                                           
 
                tmr_registers(0)(838)    <= not(local_tmr_voter(837));                                                                           
                tmr_registers(1)(838)    <= not(local_tmr_voter(837));                                                                           
                tmr_registers(2)(838)    <= not(local_tmr_voter(837));                                                                           
 
                tmr_registers(0)(839)    <= not(local_tmr_voter(838));                                                                           
                tmr_registers(1)(839)    <= not(local_tmr_voter(838));                                                                           
                tmr_registers(2)(839)    <= not(local_tmr_voter(838));                                                                           
 
                tmr_registers(0)(840)    <= not(local_tmr_voter(839));                                                                           
                tmr_registers(1)(840)    <= not(local_tmr_voter(839));                                                                           
                tmr_registers(2)(840)    <= not(local_tmr_voter(839));                                                                           
 
                tmr_registers(0)(841)    <= not(local_tmr_voter(840));                                                                           
                tmr_registers(1)(841)    <= not(local_tmr_voter(840));                                                                           
                tmr_registers(2)(841)    <= not(local_tmr_voter(840));                                                                           
 
                tmr_registers(0)(842)    <= not(local_tmr_voter(841));                                                                           
                tmr_registers(1)(842)    <= not(local_tmr_voter(841));                                                                           
                tmr_registers(2)(842)    <= not(local_tmr_voter(841));                                                                           
 
                tmr_registers(0)(843)    <= not(local_tmr_voter(842));                                                                           
                tmr_registers(1)(843)    <= not(local_tmr_voter(842));                                                                           
                tmr_registers(2)(843)    <= not(local_tmr_voter(842));                                                                           
 
                tmr_registers(0)(844)    <= not(local_tmr_voter(843));                                                                           
                tmr_registers(1)(844)    <= not(local_tmr_voter(843));                                                                           
                tmr_registers(2)(844)    <= not(local_tmr_voter(843));                                                                           
 
                tmr_registers(0)(845)    <= not(local_tmr_voter(844));                                                                           
                tmr_registers(1)(845)    <= not(local_tmr_voter(844));                                                                           
                tmr_registers(2)(845)    <= not(local_tmr_voter(844));                                                                           
 
                tmr_registers(0)(846)    <= not(local_tmr_voter(845));                                                                           
                tmr_registers(1)(846)    <= not(local_tmr_voter(845));                                                                           
                tmr_registers(2)(846)    <= not(local_tmr_voter(845));                                                                           
 
                tmr_registers(0)(847)    <= not(local_tmr_voter(846));                                                                           
                tmr_registers(1)(847)    <= not(local_tmr_voter(846));                                                                           
                tmr_registers(2)(847)    <= not(local_tmr_voter(846));                                                                           
 
                tmr_registers(0)(848)    <= not(local_tmr_voter(847));                                                                           
                tmr_registers(1)(848)    <= not(local_tmr_voter(847));                                                                           
                tmr_registers(2)(848)    <= not(local_tmr_voter(847));                                                                           
 
                tmr_registers(0)(849)    <= not(local_tmr_voter(848));                                                                           
                tmr_registers(1)(849)    <= not(local_tmr_voter(848));                                                                           
                tmr_registers(2)(849)    <= not(local_tmr_voter(848));                                                                           
 
                tmr_registers(0)(850)    <= not(local_tmr_voter(849));                                                                           
                tmr_registers(1)(850)    <= not(local_tmr_voter(849));                                                                           
                tmr_registers(2)(850)    <= not(local_tmr_voter(849));                                                                           
 
                tmr_registers(0)(851)    <= not(local_tmr_voter(850));                                                                           
                tmr_registers(1)(851)    <= not(local_tmr_voter(850));                                                                           
                tmr_registers(2)(851)    <= not(local_tmr_voter(850));                                                                           
 
                tmr_registers(0)(852)    <= not(local_tmr_voter(851));                                                                           
                tmr_registers(1)(852)    <= not(local_tmr_voter(851));                                                                           
                tmr_registers(2)(852)    <= not(local_tmr_voter(851));                                                                           
 
                tmr_registers(0)(853)    <= not(local_tmr_voter(852));                                                                           
                tmr_registers(1)(853)    <= not(local_tmr_voter(852));                                                                           
                tmr_registers(2)(853)    <= not(local_tmr_voter(852));                                                                           
 
                tmr_registers(0)(854)    <= not(local_tmr_voter(853));                                                                           
                tmr_registers(1)(854)    <= not(local_tmr_voter(853));                                                                           
                tmr_registers(2)(854)    <= not(local_tmr_voter(853));                                                                           
 
                tmr_registers(0)(855)    <= not(local_tmr_voter(854));                                                                           
                tmr_registers(1)(855)    <= not(local_tmr_voter(854));                                                                           
                tmr_registers(2)(855)    <= not(local_tmr_voter(854));                                                                           
 
                tmr_registers(0)(856)    <= not(local_tmr_voter(855));                                                                           
                tmr_registers(1)(856)    <= not(local_tmr_voter(855));                                                                           
                tmr_registers(2)(856)    <= not(local_tmr_voter(855));                                                                           
 
                tmr_registers(0)(857)    <= not(local_tmr_voter(856));                                                                           
                tmr_registers(1)(857)    <= not(local_tmr_voter(856));                                                                           
                tmr_registers(2)(857)    <= not(local_tmr_voter(856));                                                                           
 
                tmr_registers(0)(858)    <= not(local_tmr_voter(857));                                                                           
                tmr_registers(1)(858)    <= not(local_tmr_voter(857));                                                                           
                tmr_registers(2)(858)    <= not(local_tmr_voter(857));                                                                           
 
                tmr_registers(0)(859)    <= not(local_tmr_voter(858));                                                                           
                tmr_registers(1)(859)    <= not(local_tmr_voter(858));                                                                           
                tmr_registers(2)(859)    <= not(local_tmr_voter(858));                                                                           
 
                tmr_registers(0)(860)    <= not(local_tmr_voter(859));                                                                           
                tmr_registers(1)(860)    <= not(local_tmr_voter(859));                                                                           
                tmr_registers(2)(860)    <= not(local_tmr_voter(859));                                                                           
 
                tmr_registers(0)(861)    <= not(local_tmr_voter(860));                                                                           
                tmr_registers(1)(861)    <= not(local_tmr_voter(860));                                                                           
                tmr_registers(2)(861)    <= not(local_tmr_voter(860));                                                                           
 
                tmr_registers(0)(862)    <= not(local_tmr_voter(861));                                                                           
                tmr_registers(1)(862)    <= not(local_tmr_voter(861));                                                                           
                tmr_registers(2)(862)    <= not(local_tmr_voter(861));                                                                           
 
                tmr_registers(0)(863)    <= not(local_tmr_voter(862));                                                                           
                tmr_registers(1)(863)    <= not(local_tmr_voter(862));                                                                           
                tmr_registers(2)(863)    <= not(local_tmr_voter(862));                                                                           
 
                tmr_registers(0)(864)    <= not(local_tmr_voter(863));                                                                           
                tmr_registers(1)(864)    <= not(local_tmr_voter(863));                                                                           
                tmr_registers(2)(864)    <= not(local_tmr_voter(863));                                                                           
 
                tmr_registers(0)(865)    <= not(local_tmr_voter(864));                                                                           
                tmr_registers(1)(865)    <= not(local_tmr_voter(864));                                                                           
                tmr_registers(2)(865)    <= not(local_tmr_voter(864));                                                                           
 
                tmr_registers(0)(866)    <= not(local_tmr_voter(865));                                                                           
                tmr_registers(1)(866)    <= not(local_tmr_voter(865));                                                                           
                tmr_registers(2)(866)    <= not(local_tmr_voter(865));                                                                           
 
                tmr_registers(0)(867)    <= not(local_tmr_voter(866));                                                                           
                tmr_registers(1)(867)    <= not(local_tmr_voter(866));                                                                           
                tmr_registers(2)(867)    <= not(local_tmr_voter(866));                                                                           
 
                tmr_registers(0)(868)    <= not(local_tmr_voter(867));                                                                           
                tmr_registers(1)(868)    <= not(local_tmr_voter(867));                                                                           
                tmr_registers(2)(868)    <= not(local_tmr_voter(867));                                                                           
 
                tmr_registers(0)(869)    <= not(local_tmr_voter(868));                                                                           
                tmr_registers(1)(869)    <= not(local_tmr_voter(868));                                                                           
                tmr_registers(2)(869)    <= not(local_tmr_voter(868));                                                                           
 
                tmr_registers(0)(870)    <= not(local_tmr_voter(869));                                                                           
                tmr_registers(1)(870)    <= not(local_tmr_voter(869));                                                                           
                tmr_registers(2)(870)    <= not(local_tmr_voter(869));                                                                           
 
                tmr_registers(0)(871)    <= not(local_tmr_voter(870));                                                                           
                tmr_registers(1)(871)    <= not(local_tmr_voter(870));                                                                           
                tmr_registers(2)(871)    <= not(local_tmr_voter(870));                                                                           
 
                tmr_registers(0)(872)    <= not(local_tmr_voter(871));                                                                           
                tmr_registers(1)(872)    <= not(local_tmr_voter(871));                                                                           
                tmr_registers(2)(872)    <= not(local_tmr_voter(871));                                                                           
 
                tmr_registers(0)(873)    <= not(local_tmr_voter(872));                                                                           
                tmr_registers(1)(873)    <= not(local_tmr_voter(872));                                                                           
                tmr_registers(2)(873)    <= not(local_tmr_voter(872));                                                                           
 
                tmr_registers(0)(874)    <= not(local_tmr_voter(873));                                                                           
                tmr_registers(1)(874)    <= not(local_tmr_voter(873));                                                                           
                tmr_registers(2)(874)    <= not(local_tmr_voter(873));                                                                           
 
                tmr_registers(0)(875)    <= not(local_tmr_voter(874));                                                                           
                tmr_registers(1)(875)    <= not(local_tmr_voter(874));                                                                           
                tmr_registers(2)(875)    <= not(local_tmr_voter(874));                                                                           
 
                tmr_registers(0)(876)    <= not(local_tmr_voter(875));                                                                           
                tmr_registers(1)(876)    <= not(local_tmr_voter(875));                                                                           
                tmr_registers(2)(876)    <= not(local_tmr_voter(875));                                                                           
 
                tmr_registers(0)(877)    <= not(local_tmr_voter(876));                                                                           
                tmr_registers(1)(877)    <= not(local_tmr_voter(876));                                                                           
                tmr_registers(2)(877)    <= not(local_tmr_voter(876));                                                                           
 
                tmr_registers(0)(878)    <= not(local_tmr_voter(877));                                                                           
                tmr_registers(1)(878)    <= not(local_tmr_voter(877));                                                                           
                tmr_registers(2)(878)    <= not(local_tmr_voter(877));                                                                           
 
                tmr_registers(0)(879)    <= not(local_tmr_voter(878));                                                                           
                tmr_registers(1)(879)    <= not(local_tmr_voter(878));                                                                           
                tmr_registers(2)(879)    <= not(local_tmr_voter(878));                                                                           
 
                tmr_registers(0)(880)    <= not(local_tmr_voter(879));                                                                           
                tmr_registers(1)(880)    <= not(local_tmr_voter(879));                                                                           
                tmr_registers(2)(880)    <= not(local_tmr_voter(879));                                                                           
 
                tmr_registers(0)(881)    <= not(local_tmr_voter(880));                                                                           
                tmr_registers(1)(881)    <= not(local_tmr_voter(880));                                                                           
                tmr_registers(2)(881)    <= not(local_tmr_voter(880));                                                                           
 
                tmr_registers(0)(882)    <= not(local_tmr_voter(881));                                                                           
                tmr_registers(1)(882)    <= not(local_tmr_voter(881));                                                                           
                tmr_registers(2)(882)    <= not(local_tmr_voter(881));                                                                           
 
                tmr_registers(0)(883)    <= not(local_tmr_voter(882));                                                                           
                tmr_registers(1)(883)    <= not(local_tmr_voter(882));                                                                           
                tmr_registers(2)(883)    <= not(local_tmr_voter(882));                                                                           
 
                tmr_registers(0)(884)    <= not(local_tmr_voter(883));                                                                           
                tmr_registers(1)(884)    <= not(local_tmr_voter(883));                                                                           
                tmr_registers(2)(884)    <= not(local_tmr_voter(883));                                                                           
 
                tmr_registers(0)(885)    <= not(local_tmr_voter(884));                                                                           
                tmr_registers(1)(885)    <= not(local_tmr_voter(884));                                                                           
                tmr_registers(2)(885)    <= not(local_tmr_voter(884));                                                                           
 
                tmr_registers(0)(886)    <= not(local_tmr_voter(885));                                                                           
                tmr_registers(1)(886)    <= not(local_tmr_voter(885));                                                                           
                tmr_registers(2)(886)    <= not(local_tmr_voter(885));                                                                           
 
                tmr_registers(0)(887)    <= not(local_tmr_voter(886));                                                                           
                tmr_registers(1)(887)    <= not(local_tmr_voter(886));                                                                           
                tmr_registers(2)(887)    <= not(local_tmr_voter(886));                                                                           
 
                tmr_registers(0)(888)    <= not(local_tmr_voter(887));                                                                           
                tmr_registers(1)(888)    <= not(local_tmr_voter(887));                                                                           
                tmr_registers(2)(888)    <= not(local_tmr_voter(887));                                                                           
 
                tmr_registers(0)(889)    <= not(local_tmr_voter(888));                                                                           
                tmr_registers(1)(889)    <= not(local_tmr_voter(888));                                                                           
                tmr_registers(2)(889)    <= not(local_tmr_voter(888));                                                                           
 
                tmr_registers(0)(890)    <= not(local_tmr_voter(889));                                                                           
                tmr_registers(1)(890)    <= not(local_tmr_voter(889));                                                                           
                tmr_registers(2)(890)    <= not(local_tmr_voter(889));                                                                           
 
                tmr_registers(0)(891)    <= not(local_tmr_voter(890));                                                                           
                tmr_registers(1)(891)    <= not(local_tmr_voter(890));                                                                           
                tmr_registers(2)(891)    <= not(local_tmr_voter(890));                                                                           
 
                tmr_registers(0)(892)    <= not(local_tmr_voter(891));                                                                           
                tmr_registers(1)(892)    <= not(local_tmr_voter(891));                                                                           
                tmr_registers(2)(892)    <= not(local_tmr_voter(891));                                                                           
 
                tmr_registers(0)(893)    <= not(local_tmr_voter(892));                                                                           
                tmr_registers(1)(893)    <= not(local_tmr_voter(892));                                                                           
                tmr_registers(2)(893)    <= not(local_tmr_voter(892));                                                                           
 
                tmr_registers(0)(894)    <= not(local_tmr_voter(893));                                                                           
                tmr_registers(1)(894)    <= not(local_tmr_voter(893));                                                                           
                tmr_registers(2)(894)    <= not(local_tmr_voter(893));                                                                           
 
                tmr_registers(0)(895)    <= not(local_tmr_voter(894));                                                                           
                tmr_registers(1)(895)    <= not(local_tmr_voter(894));                                                                           
                tmr_registers(2)(895)    <= not(local_tmr_voter(894));                                                                           
 
                tmr_registers(0)(896)    <= not(local_tmr_voter(895));                                                                           
                tmr_registers(1)(896)    <= not(local_tmr_voter(895));                                                                           
                tmr_registers(2)(896)    <= not(local_tmr_voter(895));                                                                           
 
                tmr_registers(0)(897)    <= not(local_tmr_voter(896));                                                                           
                tmr_registers(1)(897)    <= not(local_tmr_voter(896));                                                                           
                tmr_registers(2)(897)    <= not(local_tmr_voter(896));                                                                           
 
                tmr_registers(0)(898)    <= not(local_tmr_voter(897));                                                                           
                tmr_registers(1)(898)    <= not(local_tmr_voter(897));                                                                           
                tmr_registers(2)(898)    <= not(local_tmr_voter(897));                                                                           
 
                tmr_registers(0)(899)    <= not(local_tmr_voter(898));                                                                           
                tmr_registers(1)(899)    <= not(local_tmr_voter(898));                                                                           
                tmr_registers(2)(899)    <= not(local_tmr_voter(898));                                                                           
 
                tmr_registers(0)(900)    <= not(local_tmr_voter(899));                                                                           
                tmr_registers(1)(900)    <= not(local_tmr_voter(899));                                                                           
                tmr_registers(2)(900)    <= not(local_tmr_voter(899));                                                                           
 
                tmr_registers(0)(901)    <= not(local_tmr_voter(900));                                                                           
                tmr_registers(1)(901)    <= not(local_tmr_voter(900));                                                                           
                tmr_registers(2)(901)    <= not(local_tmr_voter(900));                                                                           
 
                tmr_registers(0)(902)    <= not(local_tmr_voter(901));                                                                           
                tmr_registers(1)(902)    <= not(local_tmr_voter(901));                                                                           
                tmr_registers(2)(902)    <= not(local_tmr_voter(901));                                                                           
 
                tmr_registers(0)(903)    <= not(local_tmr_voter(902));                                                                           
                tmr_registers(1)(903)    <= not(local_tmr_voter(902));                                                                           
                tmr_registers(2)(903)    <= not(local_tmr_voter(902));                                                                           
 
                tmr_registers(0)(904)    <= not(local_tmr_voter(903));                                                                           
                tmr_registers(1)(904)    <= not(local_tmr_voter(903));                                                                           
                tmr_registers(2)(904)    <= not(local_tmr_voter(903));                                                                           
 
                tmr_registers(0)(905)    <= not(local_tmr_voter(904));                                                                           
                tmr_registers(1)(905)    <= not(local_tmr_voter(904));                                                                           
                tmr_registers(2)(905)    <= not(local_tmr_voter(904));                                                                           
 
                tmr_registers(0)(906)    <= not(local_tmr_voter(905));                                                                           
                tmr_registers(1)(906)    <= not(local_tmr_voter(905));                                                                           
                tmr_registers(2)(906)    <= not(local_tmr_voter(905));                                                                           
 
                tmr_registers(0)(907)    <= not(local_tmr_voter(906));                                                                           
                tmr_registers(1)(907)    <= not(local_tmr_voter(906));                                                                           
                tmr_registers(2)(907)    <= not(local_tmr_voter(906));                                                                           
 
                tmr_registers(0)(908)    <= not(local_tmr_voter(907));                                                                           
                tmr_registers(1)(908)    <= not(local_tmr_voter(907));                                                                           
                tmr_registers(2)(908)    <= not(local_tmr_voter(907));                                                                           
 
                tmr_registers(0)(909)    <= not(local_tmr_voter(908));                                                                           
                tmr_registers(1)(909)    <= not(local_tmr_voter(908));                                                                           
                tmr_registers(2)(909)    <= not(local_tmr_voter(908));                                                                           
 
                tmr_registers(0)(910)    <= not(local_tmr_voter(909));                                                                           
                tmr_registers(1)(910)    <= not(local_tmr_voter(909));                                                                           
                tmr_registers(2)(910)    <= not(local_tmr_voter(909));                                                                           
 
                tmr_registers(0)(911)    <= not(local_tmr_voter(910));                                                                           
                tmr_registers(1)(911)    <= not(local_tmr_voter(910));                                                                           
                tmr_registers(2)(911)    <= not(local_tmr_voter(910));                                                                           
 
                tmr_registers(0)(912)    <= not(local_tmr_voter(911));                                                                           
                tmr_registers(1)(912)    <= not(local_tmr_voter(911));                                                                           
                tmr_registers(2)(912)    <= not(local_tmr_voter(911));                                                                           
 
                tmr_registers(0)(913)    <= not(local_tmr_voter(912));                                                                           
                tmr_registers(1)(913)    <= not(local_tmr_voter(912));                                                                           
                tmr_registers(2)(913)    <= not(local_tmr_voter(912));                                                                           
 
                tmr_registers(0)(914)    <= not(local_tmr_voter(913));                                                                           
                tmr_registers(1)(914)    <= not(local_tmr_voter(913));                                                                           
                tmr_registers(2)(914)    <= not(local_tmr_voter(913));                                                                           
 
                tmr_registers(0)(915)    <= not(local_tmr_voter(914));                                                                           
                tmr_registers(1)(915)    <= not(local_tmr_voter(914));                                                                           
                tmr_registers(2)(915)    <= not(local_tmr_voter(914));                                                                           
 
                tmr_registers(0)(916)    <= not(local_tmr_voter(915));                                                                           
                tmr_registers(1)(916)    <= not(local_tmr_voter(915));                                                                           
                tmr_registers(2)(916)    <= not(local_tmr_voter(915));                                                                           
 
                tmr_registers(0)(917)    <= not(local_tmr_voter(916));                                                                           
                tmr_registers(1)(917)    <= not(local_tmr_voter(916));                                                                           
                tmr_registers(2)(917)    <= not(local_tmr_voter(916));                                                                           
 
                tmr_registers(0)(918)    <= not(local_tmr_voter(917));                                                                           
                tmr_registers(1)(918)    <= not(local_tmr_voter(917));                                                                           
                tmr_registers(2)(918)    <= not(local_tmr_voter(917));                                                                           
 
                tmr_registers(0)(919)    <= not(local_tmr_voter(918));                                                                           
                tmr_registers(1)(919)    <= not(local_tmr_voter(918));                                                                           
                tmr_registers(2)(919)    <= not(local_tmr_voter(918));                                                                           
 
                tmr_registers(0)(920)    <= not(local_tmr_voter(919));                                                                           
                tmr_registers(1)(920)    <= not(local_tmr_voter(919));                                                                           
                tmr_registers(2)(920)    <= not(local_tmr_voter(919));                                                                           
 
                tmr_registers(0)(921)    <= not(local_tmr_voter(920));                                                                           
                tmr_registers(1)(921)    <= not(local_tmr_voter(920));                                                                           
                tmr_registers(2)(921)    <= not(local_tmr_voter(920));                                                                           
 
                tmr_registers(0)(922)    <= not(local_tmr_voter(921));                                                                           
                tmr_registers(1)(922)    <= not(local_tmr_voter(921));                                                                           
                tmr_registers(2)(922)    <= not(local_tmr_voter(921));                                                                           
 
                tmr_registers(0)(923)    <= not(local_tmr_voter(922));                                                                           
                tmr_registers(1)(923)    <= not(local_tmr_voter(922));                                                                           
                tmr_registers(2)(923)    <= not(local_tmr_voter(922));                                                                           
 
                tmr_registers(0)(924)    <= not(local_tmr_voter(923));                                                                           
                tmr_registers(1)(924)    <= not(local_tmr_voter(923));                                                                           
                tmr_registers(2)(924)    <= not(local_tmr_voter(923));                                                                           
 
                tmr_registers(0)(925)    <= not(local_tmr_voter(924));                                                                           
                tmr_registers(1)(925)    <= not(local_tmr_voter(924));                                                                           
                tmr_registers(2)(925)    <= not(local_tmr_voter(924));                                                                           
 
                tmr_registers(0)(926)    <= not(local_tmr_voter(925));                                                                           
                tmr_registers(1)(926)    <= not(local_tmr_voter(925));                                                                           
                tmr_registers(2)(926)    <= not(local_tmr_voter(925));                                                                           
 
                tmr_registers(0)(927)    <= not(local_tmr_voter(926));                                                                           
                tmr_registers(1)(927)    <= not(local_tmr_voter(926));                                                                           
                tmr_registers(2)(927)    <= not(local_tmr_voter(926));                                                                           
 
                tmr_registers(0)(928)    <= not(local_tmr_voter(927));                                                                           
                tmr_registers(1)(928)    <= not(local_tmr_voter(927));                                                                           
                tmr_registers(2)(928)    <= not(local_tmr_voter(927));                                                                           
 
                tmr_registers(0)(929)    <= not(local_tmr_voter(928));                                                                           
                tmr_registers(1)(929)    <= not(local_tmr_voter(928));                                                                           
                tmr_registers(2)(929)    <= not(local_tmr_voter(928));                                                                           
 
                tmr_registers(0)(930)    <= not(local_tmr_voter(929));                                                                           
                tmr_registers(1)(930)    <= not(local_tmr_voter(929));                                                                           
                tmr_registers(2)(930)    <= not(local_tmr_voter(929));                                                                           
 
                tmr_registers(0)(931)    <= not(local_tmr_voter(930));                                                                           
                tmr_registers(1)(931)    <= not(local_tmr_voter(930));                                                                           
                tmr_registers(2)(931)    <= not(local_tmr_voter(930));                                                                           
 
                tmr_registers(0)(932)    <= not(local_tmr_voter(931));                                                                           
                tmr_registers(1)(932)    <= not(local_tmr_voter(931));                                                                           
                tmr_registers(2)(932)    <= not(local_tmr_voter(931));                                                                           
 
                tmr_registers(0)(933)    <= not(local_tmr_voter(932));                                                                           
                tmr_registers(1)(933)    <= not(local_tmr_voter(932));                                                                           
                tmr_registers(2)(933)    <= not(local_tmr_voter(932));                                                                           
 
                tmr_registers(0)(934)    <= not(local_tmr_voter(933));                                                                           
                tmr_registers(1)(934)    <= not(local_tmr_voter(933));                                                                           
                tmr_registers(2)(934)    <= not(local_tmr_voter(933));                                                                           
 
                tmr_registers(0)(935)    <= not(local_tmr_voter(934));                                                                           
                tmr_registers(1)(935)    <= not(local_tmr_voter(934));                                                                           
                tmr_registers(2)(935)    <= not(local_tmr_voter(934));                                                                           
 
                tmr_registers(0)(936)    <= not(local_tmr_voter(935));                                                                           
                tmr_registers(1)(936)    <= not(local_tmr_voter(935));                                                                           
                tmr_registers(2)(936)    <= not(local_tmr_voter(935));                                                                           
 
                tmr_registers(0)(937)    <= not(local_tmr_voter(936));                                                                           
                tmr_registers(1)(937)    <= not(local_tmr_voter(936));                                                                           
                tmr_registers(2)(937)    <= not(local_tmr_voter(936));                                                                           
 
                tmr_registers(0)(938)    <= not(local_tmr_voter(937));                                                                           
                tmr_registers(1)(938)    <= not(local_tmr_voter(937));                                                                           
                tmr_registers(2)(938)    <= not(local_tmr_voter(937));                                                                           
 
                tmr_registers(0)(939)    <= not(local_tmr_voter(938));                                                                           
                tmr_registers(1)(939)    <= not(local_tmr_voter(938));                                                                           
                tmr_registers(2)(939)    <= not(local_tmr_voter(938));                                                                           
 
                tmr_registers(0)(940)    <= not(local_tmr_voter(939));                                                                           
                tmr_registers(1)(940)    <= not(local_tmr_voter(939));                                                                           
                tmr_registers(2)(940)    <= not(local_tmr_voter(939));                                                                           
 
                tmr_registers(0)(941)    <= not(local_tmr_voter(940));                                                                           
                tmr_registers(1)(941)    <= not(local_tmr_voter(940));                                                                           
                tmr_registers(2)(941)    <= not(local_tmr_voter(940));                                                                           
 
                tmr_registers(0)(942)    <= not(local_tmr_voter(941));                                                                           
                tmr_registers(1)(942)    <= not(local_tmr_voter(941));                                                                           
                tmr_registers(2)(942)    <= not(local_tmr_voter(941));                                                                           
 
                tmr_registers(0)(943)    <= not(local_tmr_voter(942));                                                                           
                tmr_registers(1)(943)    <= not(local_tmr_voter(942));                                                                           
                tmr_registers(2)(943)    <= not(local_tmr_voter(942));                                                                           
 
                tmr_registers(0)(944)    <= not(local_tmr_voter(943));                                                                           
                tmr_registers(1)(944)    <= not(local_tmr_voter(943));                                                                           
                tmr_registers(2)(944)    <= not(local_tmr_voter(943));                                                                           
 
                tmr_registers(0)(945)    <= not(local_tmr_voter(944));                                                                           
                tmr_registers(1)(945)    <= not(local_tmr_voter(944));                                                                           
                tmr_registers(2)(945)    <= not(local_tmr_voter(944));                                                                           
 
                tmr_registers(0)(946)    <= not(local_tmr_voter(945));                                                                           
                tmr_registers(1)(946)    <= not(local_tmr_voter(945));                                                                           
                tmr_registers(2)(946)    <= not(local_tmr_voter(945));                                                                           
 
                tmr_registers(0)(947)    <= not(local_tmr_voter(946));                                                                           
                tmr_registers(1)(947)    <= not(local_tmr_voter(946));                                                                           
                tmr_registers(2)(947)    <= not(local_tmr_voter(946));                                                                           
 
                tmr_registers(0)(948)    <= not(local_tmr_voter(947));                                                                           
                tmr_registers(1)(948)    <= not(local_tmr_voter(947));                                                                           
                tmr_registers(2)(948)    <= not(local_tmr_voter(947));                                                                           
 
                tmr_registers(0)(949)    <= not(local_tmr_voter(948));                                                                           
                tmr_registers(1)(949)    <= not(local_tmr_voter(948));                                                                           
                tmr_registers(2)(949)    <= not(local_tmr_voter(948));                                                                           
 
                tmr_registers(0)(950)    <= not(local_tmr_voter(949));                                                                           
                tmr_registers(1)(950)    <= not(local_tmr_voter(949));                                                                           
                tmr_registers(2)(950)    <= not(local_tmr_voter(949));                                                                           
 
                tmr_registers(0)(951)    <= not(local_tmr_voter(950));                                                                           
                tmr_registers(1)(951)    <= not(local_tmr_voter(950));                                                                           
                tmr_registers(2)(951)    <= not(local_tmr_voter(950));                                                                           
 
                tmr_registers(0)(952)    <= not(local_tmr_voter(951));                                                                           
                tmr_registers(1)(952)    <= not(local_tmr_voter(951));                                                                           
                tmr_registers(2)(952)    <= not(local_tmr_voter(951));                                                                           
 
                tmr_registers(0)(953)    <= not(local_tmr_voter(952));                                                                           
                tmr_registers(1)(953)    <= not(local_tmr_voter(952));                                                                           
                tmr_registers(2)(953)    <= not(local_tmr_voter(952));                                                                           
 
                tmr_registers(0)(954)    <= not(local_tmr_voter(953));                                                                           
                tmr_registers(1)(954)    <= not(local_tmr_voter(953));                                                                           
                tmr_registers(2)(954)    <= not(local_tmr_voter(953));                                                                           
 
                tmr_registers(0)(955)    <= not(local_tmr_voter(954));                                                                           
                tmr_registers(1)(955)    <= not(local_tmr_voter(954));                                                                           
                tmr_registers(2)(955)    <= not(local_tmr_voter(954));                                                                           
 
                tmr_registers(0)(956)    <= not(local_tmr_voter(955));                                                                           
                tmr_registers(1)(956)    <= not(local_tmr_voter(955));                                                                           
                tmr_registers(2)(956)    <= not(local_tmr_voter(955));                                                                           
 
                tmr_registers(0)(957)    <= not(local_tmr_voter(956));                                                                           
                tmr_registers(1)(957)    <= not(local_tmr_voter(956));                                                                           
                tmr_registers(2)(957)    <= not(local_tmr_voter(956));                                                                           
 
                tmr_registers(0)(958)    <= not(local_tmr_voter(957));                                                                           
                tmr_registers(1)(958)    <= not(local_tmr_voter(957));                                                                           
                tmr_registers(2)(958)    <= not(local_tmr_voter(957));                                                                           
 
                tmr_registers(0)(959)    <= not(local_tmr_voter(958));                                                                           
                tmr_registers(1)(959)    <= not(local_tmr_voter(958));                                                                           
                tmr_registers(2)(959)    <= not(local_tmr_voter(958));                                                                           
 
                tmr_registers(0)(960)    <= not(local_tmr_voter(959));                                                                           
                tmr_registers(1)(960)    <= not(local_tmr_voter(959));                                                                           
                tmr_registers(2)(960)    <= not(local_tmr_voter(959));                                                                           
 
                tmr_registers(0)(961)    <= not(local_tmr_voter(960));                                                                           
                tmr_registers(1)(961)    <= not(local_tmr_voter(960));                                                                           
                tmr_registers(2)(961)    <= not(local_tmr_voter(960));                                                                           
 
                tmr_registers(0)(962)    <= not(local_tmr_voter(961));                                                                           
                tmr_registers(1)(962)    <= not(local_tmr_voter(961));                                                                           
                tmr_registers(2)(962)    <= not(local_tmr_voter(961));                                                                           
 
                tmr_registers(0)(963)    <= not(local_tmr_voter(962));                                                                           
                tmr_registers(1)(963)    <= not(local_tmr_voter(962));                                                                           
                tmr_registers(2)(963)    <= not(local_tmr_voter(962));                                                                           
 
                tmr_registers(0)(964)    <= not(local_tmr_voter(963));                                                                           
                tmr_registers(1)(964)    <= not(local_tmr_voter(963));                                                                           
                tmr_registers(2)(964)    <= not(local_tmr_voter(963));                                                                           
 
                tmr_registers(0)(965)    <= not(local_tmr_voter(964));                                                                           
                tmr_registers(1)(965)    <= not(local_tmr_voter(964));                                                                           
                tmr_registers(2)(965)    <= not(local_tmr_voter(964));                                                                           
 
                tmr_registers(0)(966)    <= not(local_tmr_voter(965));                                                                           
                tmr_registers(1)(966)    <= not(local_tmr_voter(965));                                                                           
                tmr_registers(2)(966)    <= not(local_tmr_voter(965));                                                                           
 
                tmr_registers(0)(967)    <= not(local_tmr_voter(966));                                                                           
                tmr_registers(1)(967)    <= not(local_tmr_voter(966));                                                                           
                tmr_registers(2)(967)    <= not(local_tmr_voter(966));                                                                           
 
                tmr_registers(0)(968)    <= not(local_tmr_voter(967));                                                                           
                tmr_registers(1)(968)    <= not(local_tmr_voter(967));                                                                           
                tmr_registers(2)(968)    <= not(local_tmr_voter(967));                                                                           
 
                tmr_registers(0)(969)    <= not(local_tmr_voter(968));                                                                           
                tmr_registers(1)(969)    <= not(local_tmr_voter(968));                                                                           
                tmr_registers(2)(969)    <= not(local_tmr_voter(968));                                                                           
 
                tmr_registers(0)(970)    <= not(local_tmr_voter(969));                                                                           
                tmr_registers(1)(970)    <= not(local_tmr_voter(969));                                                                           
                tmr_registers(2)(970)    <= not(local_tmr_voter(969));                                                                           
 
                tmr_registers(0)(971)    <= not(local_tmr_voter(970));                                                                           
                tmr_registers(1)(971)    <= not(local_tmr_voter(970));                                                                           
                tmr_registers(2)(971)    <= not(local_tmr_voter(970));                                                                           
 
                tmr_registers(0)(972)    <= not(local_tmr_voter(971));                                                                           
                tmr_registers(1)(972)    <= not(local_tmr_voter(971));                                                                           
                tmr_registers(2)(972)    <= not(local_tmr_voter(971));                                                                           
 
                tmr_registers(0)(973)    <= not(local_tmr_voter(972));                                                                           
                tmr_registers(1)(973)    <= not(local_tmr_voter(972));                                                                           
                tmr_registers(2)(973)    <= not(local_tmr_voter(972));                                                                           
 
                tmr_registers(0)(974)    <= not(local_tmr_voter(973));                                                                           
                tmr_registers(1)(974)    <= not(local_tmr_voter(973));                                                                           
                tmr_registers(2)(974)    <= not(local_tmr_voter(973));                                                                           
 
                tmr_registers(0)(975)    <= not(local_tmr_voter(974));                                                                           
                tmr_registers(1)(975)    <= not(local_tmr_voter(974));                                                                           
                tmr_registers(2)(975)    <= not(local_tmr_voter(974));                                                                           
 
                tmr_registers(0)(976)    <= not(local_tmr_voter(975));                                                                           
                tmr_registers(1)(976)    <= not(local_tmr_voter(975));                                                                           
                tmr_registers(2)(976)    <= not(local_tmr_voter(975));                                                                           
 
                tmr_registers(0)(977)    <= not(local_tmr_voter(976));                                                                           
                tmr_registers(1)(977)    <= not(local_tmr_voter(976));                                                                           
                tmr_registers(2)(977)    <= not(local_tmr_voter(976));                                                                           
 
                tmr_registers(0)(978)    <= not(local_tmr_voter(977));                                                                           
                tmr_registers(1)(978)    <= not(local_tmr_voter(977));                                                                           
                tmr_registers(2)(978)    <= not(local_tmr_voter(977));                                                                           
 
                tmr_registers(0)(979)    <= not(local_tmr_voter(978));                                                                           
                tmr_registers(1)(979)    <= not(local_tmr_voter(978));                                                                           
                tmr_registers(2)(979)    <= not(local_tmr_voter(978));                                                                           
 
                tmr_registers(0)(980)    <= not(local_tmr_voter(979));                                                                           
                tmr_registers(1)(980)    <= not(local_tmr_voter(979));                                                                           
                tmr_registers(2)(980)    <= not(local_tmr_voter(979));                                                                           
 
                tmr_registers(0)(981)    <= not(local_tmr_voter(980));                                                                           
                tmr_registers(1)(981)    <= not(local_tmr_voter(980));                                                                           
                tmr_registers(2)(981)    <= not(local_tmr_voter(980));                                                                           
 
                tmr_registers(0)(982)    <= not(local_tmr_voter(981));                                                                           
                tmr_registers(1)(982)    <= not(local_tmr_voter(981));                                                                           
                tmr_registers(2)(982)    <= not(local_tmr_voter(981));                                                                           
 
                tmr_registers(0)(983)    <= not(local_tmr_voter(982));                                                                           
                tmr_registers(1)(983)    <= not(local_tmr_voter(982));                                                                           
                tmr_registers(2)(983)    <= not(local_tmr_voter(982));                                                                           
 
                tmr_registers(0)(984)    <= not(local_tmr_voter(983));                                                                           
                tmr_registers(1)(984)    <= not(local_tmr_voter(983));                                                                           
                tmr_registers(2)(984)    <= not(local_tmr_voter(983));                                                                           
 
                tmr_registers(0)(985)    <= not(local_tmr_voter(984));                                                                           
                tmr_registers(1)(985)    <= not(local_tmr_voter(984));                                                                           
                tmr_registers(2)(985)    <= not(local_tmr_voter(984));                                                                           
 
                tmr_registers(0)(986)    <= not(local_tmr_voter(985));                                                                           
                tmr_registers(1)(986)    <= not(local_tmr_voter(985));                                                                           
                tmr_registers(2)(986)    <= not(local_tmr_voter(985));                                                                           
 
                tmr_registers(0)(987)    <= not(local_tmr_voter(986));                                                                           
                tmr_registers(1)(987)    <= not(local_tmr_voter(986));                                                                           
                tmr_registers(2)(987)    <= not(local_tmr_voter(986));                                                                           
 
                tmr_registers(0)(988)    <= not(local_tmr_voter(987));                                                                           
                tmr_registers(1)(988)    <= not(local_tmr_voter(987));                                                                           
                tmr_registers(2)(988)    <= not(local_tmr_voter(987));                                                                           
 
                tmr_registers(0)(989)    <= not(local_tmr_voter(988));                                                                           
                tmr_registers(1)(989)    <= not(local_tmr_voter(988));                                                                           
                tmr_registers(2)(989)    <= not(local_tmr_voter(988));                                                                           
 
                tmr_registers(0)(990)    <= not(local_tmr_voter(989));                                                                           
                tmr_registers(1)(990)    <= not(local_tmr_voter(989));                                                                           
                tmr_registers(2)(990)    <= not(local_tmr_voter(989));                                                                           
 
                tmr_registers(0)(991)    <= not(local_tmr_voter(990));                                                                           
                tmr_registers(1)(991)    <= not(local_tmr_voter(990));                                                                           
                tmr_registers(2)(991)    <= not(local_tmr_voter(990));                                                                           
 
                tmr_registers(0)(992)    <= not(local_tmr_voter(991));                                                                           
                tmr_registers(1)(992)    <= not(local_tmr_voter(991));                                                                           
                tmr_registers(2)(992)    <= not(local_tmr_voter(991));                                                                           
 
                tmr_registers(0)(993)    <= not(local_tmr_voter(992));                                                                           
                tmr_registers(1)(993)    <= not(local_tmr_voter(992));                                                                           
                tmr_registers(2)(993)    <= not(local_tmr_voter(992));                                                                           
 
                tmr_registers(0)(994)    <= not(local_tmr_voter(993));                                                                           
                tmr_registers(1)(994)    <= not(local_tmr_voter(993));                                                                           
                tmr_registers(2)(994)    <= not(local_tmr_voter(993));                                                                           
 
                tmr_registers(0)(995)    <= not(local_tmr_voter(994));                                                                           
                tmr_registers(1)(995)    <= not(local_tmr_voter(994));                                                                           
                tmr_registers(2)(995)    <= not(local_tmr_voter(994));                                                                           
 
                tmr_registers(0)(996)    <= not(local_tmr_voter(995));                                                                           
                tmr_registers(1)(996)    <= not(local_tmr_voter(995));                                                                           
                tmr_registers(2)(996)    <= not(local_tmr_voter(995));                                                                           
 
                tmr_registers(0)(997)    <= not(local_tmr_voter(996));                                                                           
                tmr_registers(1)(997)    <= not(local_tmr_voter(996));                                                                           
                tmr_registers(2)(997)    <= not(local_tmr_voter(996));                                                                           
 
                tmr_registers(0)(998)    <= not(local_tmr_voter(997));                                                                           
                tmr_registers(1)(998)    <= not(local_tmr_voter(997));                                                                           
                tmr_registers(2)(998)    <= not(local_tmr_voter(997));                                                                           
 
                tmr_registers(0)(999)    <= not(local_tmr_voter(998));                                                                           
                tmr_registers(1)(999)    <= not(local_tmr_voter(998));                                                                           
                tmr_registers(2)(999)    <= not(local_tmr_voter(998));                                                                           
 
                                                                                                                                         
        end if;                                                                                                                          
    end process;                                                                                                                         
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Voter                                                                                                                             
    ------------------------------------------                                                                                           
                                                                                                                                         
        local_tmr_voter(0)  <= data_in;                                                                                                        
                                                                                                                                         
        local_tmr_voter(1)  <=    (tmr_registers(0)(1) and tmr_registers(1)(1)) or                                                             
                            (tmr_registers(1)(1) and tmr_registers(2)(1)) or                                                             
                            (tmr_registers(0)(1) and tmr_registers(2)(1));                                                               
                                                                                                                                         
        local_tmr_voter(2)  <=    (tmr_registers(0)(2) and tmr_registers(1)(2)) or                                                             
                            (tmr_registers(1)(2) and tmr_registers(2)(2)) or                                                             
                            (tmr_registers(0)(2) and tmr_registers(2)(2));                                                               
                                                                                                                                         
        local_tmr_voter(3)  <=    (tmr_registers(0)(3) and tmr_registers(1)(3)) or                                                             
                            (tmr_registers(1)(3) and tmr_registers(2)(3)) or                                                             
                            (tmr_registers(0)(3) and tmr_registers(2)(3));                                                               
                                                                                                                                         
        local_tmr_voter(4)  <=    (tmr_registers(0)(4) and tmr_registers(1)(4)) or                                                             
                            (tmr_registers(1)(4) and tmr_registers(2)(4)) or                                                             
                            (tmr_registers(0)(4) and tmr_registers(2)(4));                                                               
                                                                                                                                         
        local_tmr_voter(5)  <=    (tmr_registers(0)(5) and tmr_registers(1)(5)) or                                                             
                            (tmr_registers(1)(5) and tmr_registers(2)(5)) or                                                             
                            (tmr_registers(0)(5) and tmr_registers(2)(5));                                                               
                                                                                                                                         
        local_tmr_voter(6)  <=    (tmr_registers(0)(6) and tmr_registers(1)(6)) or                                                             
                            (tmr_registers(1)(6) and tmr_registers(2)(6)) or                                                             
                            (tmr_registers(0)(6) and tmr_registers(2)(6));                                                               
                                                                                                                                         
        local_tmr_voter(7)  <=    (tmr_registers(0)(7) and tmr_registers(1)(7)) or                                                             
                            (tmr_registers(1)(7) and tmr_registers(2)(7)) or                                                             
                            (tmr_registers(0)(7) and tmr_registers(2)(7));                                                               
                                                                                                                                         
        local_tmr_voter(8)  <=    (tmr_registers(0)(8) and tmr_registers(1)(8)) or                                                             
                            (tmr_registers(1)(8) and tmr_registers(2)(8)) or                                                             
                            (tmr_registers(0)(8) and tmr_registers(2)(8));                                                               
                                                                                                                                         
        local_tmr_voter(9)  <=    (tmr_registers(0)(9) and tmr_registers(1)(9)) or                                                             
                            (tmr_registers(1)(9) and tmr_registers(2)(9)) or                                                             
                            (tmr_registers(0)(9) and tmr_registers(2)(9));                                                               
                                                                                                                                         
        local_tmr_voter(10)  <=    (tmr_registers(0)(10) and tmr_registers(1)(10)) or                                                             
                            (tmr_registers(1)(10) and tmr_registers(2)(10)) or                                                             
                            (tmr_registers(0)(10) and tmr_registers(2)(10));                                                               
                                                                                                                                         
        local_tmr_voter(11)  <=    (tmr_registers(0)(11) and tmr_registers(1)(11)) or                                                             
                            (tmr_registers(1)(11) and tmr_registers(2)(11)) or                                                             
                            (tmr_registers(0)(11) and tmr_registers(2)(11));                                                               
                                                                                                                                         
        local_tmr_voter(12)  <=    (tmr_registers(0)(12) and tmr_registers(1)(12)) or                                                             
                            (tmr_registers(1)(12) and tmr_registers(2)(12)) or                                                             
                            (tmr_registers(0)(12) and tmr_registers(2)(12));                                                               
                                                                                                                                         
        local_tmr_voter(13)  <=    (tmr_registers(0)(13) and tmr_registers(1)(13)) or                                                             
                            (tmr_registers(1)(13) and tmr_registers(2)(13)) or                                                             
                            (tmr_registers(0)(13) and tmr_registers(2)(13));                                                               
                                                                                                                                         
        local_tmr_voter(14)  <=    (tmr_registers(0)(14) and tmr_registers(1)(14)) or                                                             
                            (tmr_registers(1)(14) and tmr_registers(2)(14)) or                                                             
                            (tmr_registers(0)(14) and tmr_registers(2)(14));                                                               
                                                                                                                                         
        local_tmr_voter(15)  <=    (tmr_registers(0)(15) and tmr_registers(1)(15)) or                                                             
                            (tmr_registers(1)(15) and tmr_registers(2)(15)) or                                                             
                            (tmr_registers(0)(15) and tmr_registers(2)(15));                                                               
                                                                                                                                         
        local_tmr_voter(16)  <=    (tmr_registers(0)(16) and tmr_registers(1)(16)) or                                                             
                            (tmr_registers(1)(16) and tmr_registers(2)(16)) or                                                             
                            (tmr_registers(0)(16) and tmr_registers(2)(16));                                                               
                                                                                                                                         
        local_tmr_voter(17)  <=    (tmr_registers(0)(17) and tmr_registers(1)(17)) or                                                             
                            (tmr_registers(1)(17) and tmr_registers(2)(17)) or                                                             
                            (tmr_registers(0)(17) and tmr_registers(2)(17));                                                               
                                                                                                                                         
        local_tmr_voter(18)  <=    (tmr_registers(0)(18) and tmr_registers(1)(18)) or                                                             
                            (tmr_registers(1)(18) and tmr_registers(2)(18)) or                                                             
                            (tmr_registers(0)(18) and tmr_registers(2)(18));                                                               
                                                                                                                                         
        local_tmr_voter(19)  <=    (tmr_registers(0)(19) and tmr_registers(1)(19)) or                                                             
                            (tmr_registers(1)(19) and tmr_registers(2)(19)) or                                                             
                            (tmr_registers(0)(19) and tmr_registers(2)(19));                                                               
                                                                                                                                         
        local_tmr_voter(20)  <=    (tmr_registers(0)(20) and tmr_registers(1)(20)) or                                                             
                            (tmr_registers(1)(20) and tmr_registers(2)(20)) or                                                             
                            (tmr_registers(0)(20) and tmr_registers(2)(20));                                                               
                                                                                                                                         
        local_tmr_voter(21)  <=    (tmr_registers(0)(21) and tmr_registers(1)(21)) or                                                             
                            (tmr_registers(1)(21) and tmr_registers(2)(21)) or                                                             
                            (tmr_registers(0)(21) and tmr_registers(2)(21));                                                               
                                                                                                                                         
        local_tmr_voter(22)  <=    (tmr_registers(0)(22) and tmr_registers(1)(22)) or                                                             
                            (tmr_registers(1)(22) and tmr_registers(2)(22)) or                                                             
                            (tmr_registers(0)(22) and tmr_registers(2)(22));                                                               
                                                                                                                                         
        local_tmr_voter(23)  <=    (tmr_registers(0)(23) and tmr_registers(1)(23)) or                                                             
                            (tmr_registers(1)(23) and tmr_registers(2)(23)) or                                                             
                            (tmr_registers(0)(23) and tmr_registers(2)(23));                                                               
                                                                                                                                         
        local_tmr_voter(24)  <=    (tmr_registers(0)(24) and tmr_registers(1)(24)) or                                                             
                            (tmr_registers(1)(24) and tmr_registers(2)(24)) or                                                             
                            (tmr_registers(0)(24) and tmr_registers(2)(24));                                                               
                                                                                                                                         
        local_tmr_voter(25)  <=    (tmr_registers(0)(25) and tmr_registers(1)(25)) or                                                             
                            (tmr_registers(1)(25) and tmr_registers(2)(25)) or                                                             
                            (tmr_registers(0)(25) and tmr_registers(2)(25));                                                               
                                                                                                                                         
        local_tmr_voter(26)  <=    (tmr_registers(0)(26) and tmr_registers(1)(26)) or                                                             
                            (tmr_registers(1)(26) and tmr_registers(2)(26)) or                                                             
                            (tmr_registers(0)(26) and tmr_registers(2)(26));                                                               
                                                                                                                                         
        local_tmr_voter(27)  <=    (tmr_registers(0)(27) and tmr_registers(1)(27)) or                                                             
                            (tmr_registers(1)(27) and tmr_registers(2)(27)) or                                                             
                            (tmr_registers(0)(27) and tmr_registers(2)(27));                                                               
                                                                                                                                         
        local_tmr_voter(28)  <=    (tmr_registers(0)(28) and tmr_registers(1)(28)) or                                                             
                            (tmr_registers(1)(28) and tmr_registers(2)(28)) or                                                             
                            (tmr_registers(0)(28) and tmr_registers(2)(28));                                                               
                                                                                                                                         
        local_tmr_voter(29)  <=    (tmr_registers(0)(29) and tmr_registers(1)(29)) or                                                             
                            (tmr_registers(1)(29) and tmr_registers(2)(29)) or                                                             
                            (tmr_registers(0)(29) and tmr_registers(2)(29));                                                               
                                                                                                                                         
        local_tmr_voter(30)  <=    (tmr_registers(0)(30) and tmr_registers(1)(30)) or                                                             
                            (tmr_registers(1)(30) and tmr_registers(2)(30)) or                                                             
                            (tmr_registers(0)(30) and tmr_registers(2)(30));                                                               
                                                                                                                                         
        local_tmr_voter(31)  <=    (tmr_registers(0)(31) and tmr_registers(1)(31)) or                                                             
                            (tmr_registers(1)(31) and tmr_registers(2)(31)) or                                                             
                            (tmr_registers(0)(31) and tmr_registers(2)(31));                                                               
                                                                                                                                         
        local_tmr_voter(32)  <=    (tmr_registers(0)(32) and tmr_registers(1)(32)) or                                                             
                            (tmr_registers(1)(32) and tmr_registers(2)(32)) or                                                             
                            (tmr_registers(0)(32) and tmr_registers(2)(32));                                                               
                                                                                                                                         
        local_tmr_voter(33)  <=    (tmr_registers(0)(33) and tmr_registers(1)(33)) or                                                             
                            (tmr_registers(1)(33) and tmr_registers(2)(33)) or                                                             
                            (tmr_registers(0)(33) and tmr_registers(2)(33));                                                               
                                                                                                                                         
        local_tmr_voter(34)  <=    (tmr_registers(0)(34) and tmr_registers(1)(34)) or                                                             
                            (tmr_registers(1)(34) and tmr_registers(2)(34)) or                                                             
                            (tmr_registers(0)(34) and tmr_registers(2)(34));                                                               
                                                                                                                                         
        local_tmr_voter(35)  <=    (tmr_registers(0)(35) and tmr_registers(1)(35)) or                                                             
                            (tmr_registers(1)(35) and tmr_registers(2)(35)) or                                                             
                            (tmr_registers(0)(35) and tmr_registers(2)(35));                                                               
                                                                                                                                         
        local_tmr_voter(36)  <=    (tmr_registers(0)(36) and tmr_registers(1)(36)) or                                                             
                            (tmr_registers(1)(36) and tmr_registers(2)(36)) or                                                             
                            (tmr_registers(0)(36) and tmr_registers(2)(36));                                                               
                                                                                                                                         
        local_tmr_voter(37)  <=    (tmr_registers(0)(37) and tmr_registers(1)(37)) or                                                             
                            (tmr_registers(1)(37) and tmr_registers(2)(37)) or                                                             
                            (tmr_registers(0)(37) and tmr_registers(2)(37));                                                               
                                                                                                                                         
        local_tmr_voter(38)  <=    (tmr_registers(0)(38) and tmr_registers(1)(38)) or                                                             
                            (tmr_registers(1)(38) and tmr_registers(2)(38)) or                                                             
                            (tmr_registers(0)(38) and tmr_registers(2)(38));                                                               
                                                                                                                                         
        local_tmr_voter(39)  <=    (tmr_registers(0)(39) and tmr_registers(1)(39)) or                                                             
                            (tmr_registers(1)(39) and tmr_registers(2)(39)) or                                                             
                            (tmr_registers(0)(39) and tmr_registers(2)(39));                                                               
                                                                                                                                         
        local_tmr_voter(40)  <=    (tmr_registers(0)(40) and tmr_registers(1)(40)) or                                                             
                            (tmr_registers(1)(40) and tmr_registers(2)(40)) or                                                             
                            (tmr_registers(0)(40) and tmr_registers(2)(40));                                                               
                                                                                                                                         
        local_tmr_voter(41)  <=    (tmr_registers(0)(41) and tmr_registers(1)(41)) or                                                             
                            (tmr_registers(1)(41) and tmr_registers(2)(41)) or                                                             
                            (tmr_registers(0)(41) and tmr_registers(2)(41));                                                               
                                                                                                                                         
        local_tmr_voter(42)  <=    (tmr_registers(0)(42) and tmr_registers(1)(42)) or                                                             
                            (tmr_registers(1)(42) and tmr_registers(2)(42)) or                                                             
                            (tmr_registers(0)(42) and tmr_registers(2)(42));                                                               
                                                                                                                                         
        local_tmr_voter(43)  <=    (tmr_registers(0)(43) and tmr_registers(1)(43)) or                                                             
                            (tmr_registers(1)(43) and tmr_registers(2)(43)) or                                                             
                            (tmr_registers(0)(43) and tmr_registers(2)(43));                                                               
                                                                                                                                         
        local_tmr_voter(44)  <=    (tmr_registers(0)(44) and tmr_registers(1)(44)) or                                                             
                            (tmr_registers(1)(44) and tmr_registers(2)(44)) or                                                             
                            (tmr_registers(0)(44) and tmr_registers(2)(44));                                                               
                                                                                                                                         
        local_tmr_voter(45)  <=    (tmr_registers(0)(45) and tmr_registers(1)(45)) or                                                             
                            (tmr_registers(1)(45) and tmr_registers(2)(45)) or                                                             
                            (tmr_registers(0)(45) and tmr_registers(2)(45));                                                               
                                                                                                                                         
        local_tmr_voter(46)  <=    (tmr_registers(0)(46) and tmr_registers(1)(46)) or                                                             
                            (tmr_registers(1)(46) and tmr_registers(2)(46)) or                                                             
                            (tmr_registers(0)(46) and tmr_registers(2)(46));                                                               
                                                                                                                                         
        local_tmr_voter(47)  <=    (tmr_registers(0)(47) and tmr_registers(1)(47)) or                                                             
                            (tmr_registers(1)(47) and tmr_registers(2)(47)) or                                                             
                            (tmr_registers(0)(47) and tmr_registers(2)(47));                                                               
                                                                                                                                         
        local_tmr_voter(48)  <=    (tmr_registers(0)(48) and tmr_registers(1)(48)) or                                                             
                            (tmr_registers(1)(48) and tmr_registers(2)(48)) or                                                             
                            (tmr_registers(0)(48) and tmr_registers(2)(48));                                                               
                                                                                                                                         
        local_tmr_voter(49)  <=    (tmr_registers(0)(49) and tmr_registers(1)(49)) or                                                             
                            (tmr_registers(1)(49) and tmr_registers(2)(49)) or                                                             
                            (tmr_registers(0)(49) and tmr_registers(2)(49));                                                               
                                                                                                                                         
        local_tmr_voter(50)  <=    (tmr_registers(0)(50) and tmr_registers(1)(50)) or                                                             
                            (tmr_registers(1)(50) and tmr_registers(2)(50)) or                                                             
                            (tmr_registers(0)(50) and tmr_registers(2)(50));                                                               
                                                                                                                                         
        local_tmr_voter(51)  <=    (tmr_registers(0)(51) and tmr_registers(1)(51)) or                                                             
                            (tmr_registers(1)(51) and tmr_registers(2)(51)) or                                                             
                            (tmr_registers(0)(51) and tmr_registers(2)(51));                                                               
                                                                                                                                         
        local_tmr_voter(52)  <=    (tmr_registers(0)(52) and tmr_registers(1)(52)) or                                                             
                            (tmr_registers(1)(52) and tmr_registers(2)(52)) or                                                             
                            (tmr_registers(0)(52) and tmr_registers(2)(52));                                                               
                                                                                                                                         
        local_tmr_voter(53)  <=    (tmr_registers(0)(53) and tmr_registers(1)(53)) or                                                             
                            (tmr_registers(1)(53) and tmr_registers(2)(53)) or                                                             
                            (tmr_registers(0)(53) and tmr_registers(2)(53));                                                               
                                                                                                                                         
        local_tmr_voter(54)  <=    (tmr_registers(0)(54) and tmr_registers(1)(54)) or                                                             
                            (tmr_registers(1)(54) and tmr_registers(2)(54)) or                                                             
                            (tmr_registers(0)(54) and tmr_registers(2)(54));                                                               
                                                                                                                                         
        local_tmr_voter(55)  <=    (tmr_registers(0)(55) and tmr_registers(1)(55)) or                                                             
                            (tmr_registers(1)(55) and tmr_registers(2)(55)) or                                                             
                            (tmr_registers(0)(55) and tmr_registers(2)(55));                                                               
                                                                                                                                         
        local_tmr_voter(56)  <=    (tmr_registers(0)(56) and tmr_registers(1)(56)) or                                                             
                            (tmr_registers(1)(56) and tmr_registers(2)(56)) or                                                             
                            (tmr_registers(0)(56) and tmr_registers(2)(56));                                                               
                                                                                                                                         
        local_tmr_voter(57)  <=    (tmr_registers(0)(57) and tmr_registers(1)(57)) or                                                             
                            (tmr_registers(1)(57) and tmr_registers(2)(57)) or                                                             
                            (tmr_registers(0)(57) and tmr_registers(2)(57));                                                               
                                                                                                                                         
        local_tmr_voter(58)  <=    (tmr_registers(0)(58) and tmr_registers(1)(58)) or                                                             
                            (tmr_registers(1)(58) and tmr_registers(2)(58)) or                                                             
                            (tmr_registers(0)(58) and tmr_registers(2)(58));                                                               
                                                                                                                                         
        local_tmr_voter(59)  <=    (tmr_registers(0)(59) and tmr_registers(1)(59)) or                                                             
                            (tmr_registers(1)(59) and tmr_registers(2)(59)) or                                                             
                            (tmr_registers(0)(59) and tmr_registers(2)(59));                                                               
                                                                                                                                         
        local_tmr_voter(60)  <=    (tmr_registers(0)(60) and tmr_registers(1)(60)) or                                                             
                            (tmr_registers(1)(60) and tmr_registers(2)(60)) or                                                             
                            (tmr_registers(0)(60) and tmr_registers(2)(60));                                                               
                                                                                                                                         
        local_tmr_voter(61)  <=    (tmr_registers(0)(61) and tmr_registers(1)(61)) or                                                             
                            (tmr_registers(1)(61) and tmr_registers(2)(61)) or                                                             
                            (tmr_registers(0)(61) and tmr_registers(2)(61));                                                               
                                                                                                                                         
        local_tmr_voter(62)  <=    (tmr_registers(0)(62) and tmr_registers(1)(62)) or                                                             
                            (tmr_registers(1)(62) and tmr_registers(2)(62)) or                                                             
                            (tmr_registers(0)(62) and tmr_registers(2)(62));                                                               
                                                                                                                                         
        local_tmr_voter(63)  <=    (tmr_registers(0)(63) and tmr_registers(1)(63)) or                                                             
                            (tmr_registers(1)(63) and tmr_registers(2)(63)) or                                                             
                            (tmr_registers(0)(63) and tmr_registers(2)(63));                                                               
                                                                                                                                         
        local_tmr_voter(64)  <=    (tmr_registers(0)(64) and tmr_registers(1)(64)) or                                                             
                            (tmr_registers(1)(64) and tmr_registers(2)(64)) or                                                             
                            (tmr_registers(0)(64) and tmr_registers(2)(64));                                                               
                                                                                                                                         
        local_tmr_voter(65)  <=    (tmr_registers(0)(65) and tmr_registers(1)(65)) or                                                             
                            (tmr_registers(1)(65) and tmr_registers(2)(65)) or                                                             
                            (tmr_registers(0)(65) and tmr_registers(2)(65));                                                               
                                                                                                                                         
        local_tmr_voter(66)  <=    (tmr_registers(0)(66) and tmr_registers(1)(66)) or                                                             
                            (tmr_registers(1)(66) and tmr_registers(2)(66)) or                                                             
                            (tmr_registers(0)(66) and tmr_registers(2)(66));                                                               
                                                                                                                                         
        local_tmr_voter(67)  <=    (tmr_registers(0)(67) and tmr_registers(1)(67)) or                                                             
                            (tmr_registers(1)(67) and tmr_registers(2)(67)) or                                                             
                            (tmr_registers(0)(67) and tmr_registers(2)(67));                                                               
                                                                                                                                         
        local_tmr_voter(68)  <=    (tmr_registers(0)(68) and tmr_registers(1)(68)) or                                                             
                            (tmr_registers(1)(68) and tmr_registers(2)(68)) or                                                             
                            (tmr_registers(0)(68) and tmr_registers(2)(68));                                                               
                                                                                                                                         
        local_tmr_voter(69)  <=    (tmr_registers(0)(69) and tmr_registers(1)(69)) or                                                             
                            (tmr_registers(1)(69) and tmr_registers(2)(69)) or                                                             
                            (tmr_registers(0)(69) and tmr_registers(2)(69));                                                               
                                                                                                                                         
        local_tmr_voter(70)  <=    (tmr_registers(0)(70) and tmr_registers(1)(70)) or                                                             
                            (tmr_registers(1)(70) and tmr_registers(2)(70)) or                                                             
                            (tmr_registers(0)(70) and tmr_registers(2)(70));                                                               
                                                                                                                                         
        local_tmr_voter(71)  <=    (tmr_registers(0)(71) and tmr_registers(1)(71)) or                                                             
                            (tmr_registers(1)(71) and tmr_registers(2)(71)) or                                                             
                            (tmr_registers(0)(71) and tmr_registers(2)(71));                                                               
                                                                                                                                         
        local_tmr_voter(72)  <=    (tmr_registers(0)(72) and tmr_registers(1)(72)) or                                                             
                            (tmr_registers(1)(72) and tmr_registers(2)(72)) or                                                             
                            (tmr_registers(0)(72) and tmr_registers(2)(72));                                                               
                                                                                                                                         
        local_tmr_voter(73)  <=    (tmr_registers(0)(73) and tmr_registers(1)(73)) or                                                             
                            (tmr_registers(1)(73) and tmr_registers(2)(73)) or                                                             
                            (tmr_registers(0)(73) and tmr_registers(2)(73));                                                               
                                                                                                                                         
        local_tmr_voter(74)  <=    (tmr_registers(0)(74) and tmr_registers(1)(74)) or                                                             
                            (tmr_registers(1)(74) and tmr_registers(2)(74)) or                                                             
                            (tmr_registers(0)(74) and tmr_registers(2)(74));                                                               
                                                                                                                                         
        local_tmr_voter(75)  <=    (tmr_registers(0)(75) and tmr_registers(1)(75)) or                                                             
                            (tmr_registers(1)(75) and tmr_registers(2)(75)) or                                                             
                            (tmr_registers(0)(75) and tmr_registers(2)(75));                                                               
                                                                                                                                         
        local_tmr_voter(76)  <=    (tmr_registers(0)(76) and tmr_registers(1)(76)) or                                                             
                            (tmr_registers(1)(76) and tmr_registers(2)(76)) or                                                             
                            (tmr_registers(0)(76) and tmr_registers(2)(76));                                                               
                                                                                                                                         
        local_tmr_voter(77)  <=    (tmr_registers(0)(77) and tmr_registers(1)(77)) or                                                             
                            (tmr_registers(1)(77) and tmr_registers(2)(77)) or                                                             
                            (tmr_registers(0)(77) and tmr_registers(2)(77));                                                               
                                                                                                                                         
        local_tmr_voter(78)  <=    (tmr_registers(0)(78) and tmr_registers(1)(78)) or                                                             
                            (tmr_registers(1)(78) and tmr_registers(2)(78)) or                                                             
                            (tmr_registers(0)(78) and tmr_registers(2)(78));                                                               
                                                                                                                                         
        local_tmr_voter(79)  <=    (tmr_registers(0)(79) and tmr_registers(1)(79)) or                                                             
                            (tmr_registers(1)(79) and tmr_registers(2)(79)) or                                                             
                            (tmr_registers(0)(79) and tmr_registers(2)(79));                                                               
                                                                                                                                         
        local_tmr_voter(80)  <=    (tmr_registers(0)(80) and tmr_registers(1)(80)) or                                                             
                            (tmr_registers(1)(80) and tmr_registers(2)(80)) or                                                             
                            (tmr_registers(0)(80) and tmr_registers(2)(80));                                                               
                                                                                                                                         
        local_tmr_voter(81)  <=    (tmr_registers(0)(81) and tmr_registers(1)(81)) or                                                             
                            (tmr_registers(1)(81) and tmr_registers(2)(81)) or                                                             
                            (tmr_registers(0)(81) and tmr_registers(2)(81));                                                               
                                                                                                                                         
        local_tmr_voter(82)  <=    (tmr_registers(0)(82) and tmr_registers(1)(82)) or                                                             
                            (tmr_registers(1)(82) and tmr_registers(2)(82)) or                                                             
                            (tmr_registers(0)(82) and tmr_registers(2)(82));                                                               
                                                                                                                                         
        local_tmr_voter(83)  <=    (tmr_registers(0)(83) and tmr_registers(1)(83)) or                                                             
                            (tmr_registers(1)(83) and tmr_registers(2)(83)) or                                                             
                            (tmr_registers(0)(83) and tmr_registers(2)(83));                                                               
                                                                                                                                         
        local_tmr_voter(84)  <=    (tmr_registers(0)(84) and tmr_registers(1)(84)) or                                                             
                            (tmr_registers(1)(84) and tmr_registers(2)(84)) or                                                             
                            (tmr_registers(0)(84) and tmr_registers(2)(84));                                                               
                                                                                                                                         
        local_tmr_voter(85)  <=    (tmr_registers(0)(85) and tmr_registers(1)(85)) or                                                             
                            (tmr_registers(1)(85) and tmr_registers(2)(85)) or                                                             
                            (tmr_registers(0)(85) and tmr_registers(2)(85));                                                               
                                                                                                                                         
        local_tmr_voter(86)  <=    (tmr_registers(0)(86) and tmr_registers(1)(86)) or                                                             
                            (tmr_registers(1)(86) and tmr_registers(2)(86)) or                                                             
                            (tmr_registers(0)(86) and tmr_registers(2)(86));                                                               
                                                                                                                                         
        local_tmr_voter(87)  <=    (tmr_registers(0)(87) and tmr_registers(1)(87)) or                                                             
                            (tmr_registers(1)(87) and tmr_registers(2)(87)) or                                                             
                            (tmr_registers(0)(87) and tmr_registers(2)(87));                                                               
                                                                                                                                         
        local_tmr_voter(88)  <=    (tmr_registers(0)(88) and tmr_registers(1)(88)) or                                                             
                            (tmr_registers(1)(88) and tmr_registers(2)(88)) or                                                             
                            (tmr_registers(0)(88) and tmr_registers(2)(88));                                                               
                                                                                                                                         
        local_tmr_voter(89)  <=    (tmr_registers(0)(89) and tmr_registers(1)(89)) or                                                             
                            (tmr_registers(1)(89) and tmr_registers(2)(89)) or                                                             
                            (tmr_registers(0)(89) and tmr_registers(2)(89));                                                               
                                                                                                                                         
        local_tmr_voter(90)  <=    (tmr_registers(0)(90) and tmr_registers(1)(90)) or                                                             
                            (tmr_registers(1)(90) and tmr_registers(2)(90)) or                                                             
                            (tmr_registers(0)(90) and tmr_registers(2)(90));                                                               
                                                                                                                                         
        local_tmr_voter(91)  <=    (tmr_registers(0)(91) and tmr_registers(1)(91)) or                                                             
                            (tmr_registers(1)(91) and tmr_registers(2)(91)) or                                                             
                            (tmr_registers(0)(91) and tmr_registers(2)(91));                                                               
                                                                                                                                         
        local_tmr_voter(92)  <=    (tmr_registers(0)(92) and tmr_registers(1)(92)) or                                                             
                            (tmr_registers(1)(92) and tmr_registers(2)(92)) or                                                             
                            (tmr_registers(0)(92) and tmr_registers(2)(92));                                                               
                                                                                                                                         
        local_tmr_voter(93)  <=    (tmr_registers(0)(93) and tmr_registers(1)(93)) or                                                             
                            (tmr_registers(1)(93) and tmr_registers(2)(93)) or                                                             
                            (tmr_registers(0)(93) and tmr_registers(2)(93));                                                               
                                                                                                                                         
        local_tmr_voter(94)  <=    (tmr_registers(0)(94) and tmr_registers(1)(94)) or                                                             
                            (tmr_registers(1)(94) and tmr_registers(2)(94)) or                                                             
                            (tmr_registers(0)(94) and tmr_registers(2)(94));                                                               
                                                                                                                                         
        local_tmr_voter(95)  <=    (tmr_registers(0)(95) and tmr_registers(1)(95)) or                                                             
                            (tmr_registers(1)(95) and tmr_registers(2)(95)) or                                                             
                            (tmr_registers(0)(95) and tmr_registers(2)(95));                                                               
                                                                                                                                         
        local_tmr_voter(96)  <=    (tmr_registers(0)(96) and tmr_registers(1)(96)) or                                                             
                            (tmr_registers(1)(96) and tmr_registers(2)(96)) or                                                             
                            (tmr_registers(0)(96) and tmr_registers(2)(96));                                                               
                                                                                                                                         
        local_tmr_voter(97)  <=    (tmr_registers(0)(97) and tmr_registers(1)(97)) or                                                             
                            (tmr_registers(1)(97) and tmr_registers(2)(97)) or                                                             
                            (tmr_registers(0)(97) and tmr_registers(2)(97));                                                               
                                                                                                                                         
        local_tmr_voter(98)  <=    (tmr_registers(0)(98) and tmr_registers(1)(98)) or                                                             
                            (tmr_registers(1)(98) and tmr_registers(2)(98)) or                                                             
                            (tmr_registers(0)(98) and tmr_registers(2)(98));                                                               
                                                                                                                                         
        local_tmr_voter(99)  <=    (tmr_registers(0)(99) and tmr_registers(1)(99)) or                                                             
                            (tmr_registers(1)(99) and tmr_registers(2)(99)) or                                                             
                            (tmr_registers(0)(99) and tmr_registers(2)(99));                                                               
                                                                                                                                         
        local_tmr_voter(100)  <=    (tmr_registers(0)(100) and tmr_registers(1)(100)) or                                                             
                            (tmr_registers(1)(100) and tmr_registers(2)(100)) or                                                             
                            (tmr_registers(0)(100) and tmr_registers(2)(100));                                                               
                                                                                                                                         
        local_tmr_voter(101)  <=    (tmr_registers(0)(101) and tmr_registers(1)(101)) or                                                             
                            (tmr_registers(1)(101) and tmr_registers(2)(101)) or                                                             
                            (tmr_registers(0)(101) and tmr_registers(2)(101));                                                               
                                                                                                                                         
        local_tmr_voter(102)  <=    (tmr_registers(0)(102) and tmr_registers(1)(102)) or                                                             
                            (tmr_registers(1)(102) and tmr_registers(2)(102)) or                                                             
                            (tmr_registers(0)(102) and tmr_registers(2)(102));                                                               
                                                                                                                                         
        local_tmr_voter(103)  <=    (tmr_registers(0)(103) and tmr_registers(1)(103)) or                                                             
                            (tmr_registers(1)(103) and tmr_registers(2)(103)) or                                                             
                            (tmr_registers(0)(103) and tmr_registers(2)(103));                                                               
                                                                                                                                         
        local_tmr_voter(104)  <=    (tmr_registers(0)(104) and tmr_registers(1)(104)) or                                                             
                            (tmr_registers(1)(104) and tmr_registers(2)(104)) or                                                             
                            (tmr_registers(0)(104) and tmr_registers(2)(104));                                                               
                                                                                                                                         
        local_tmr_voter(105)  <=    (tmr_registers(0)(105) and tmr_registers(1)(105)) or                                                             
                            (tmr_registers(1)(105) and tmr_registers(2)(105)) or                                                             
                            (tmr_registers(0)(105) and tmr_registers(2)(105));                                                               
                                                                                                                                         
        local_tmr_voter(106)  <=    (tmr_registers(0)(106) and tmr_registers(1)(106)) or                                                             
                            (tmr_registers(1)(106) and tmr_registers(2)(106)) or                                                             
                            (tmr_registers(0)(106) and tmr_registers(2)(106));                                                               
                                                                                                                                         
        local_tmr_voter(107)  <=    (tmr_registers(0)(107) and tmr_registers(1)(107)) or                                                             
                            (tmr_registers(1)(107) and tmr_registers(2)(107)) or                                                             
                            (tmr_registers(0)(107) and tmr_registers(2)(107));                                                               
                                                                                                                                         
        local_tmr_voter(108)  <=    (tmr_registers(0)(108) and tmr_registers(1)(108)) or                                                             
                            (tmr_registers(1)(108) and tmr_registers(2)(108)) or                                                             
                            (tmr_registers(0)(108) and tmr_registers(2)(108));                                                               
                                                                                                                                         
        local_tmr_voter(109)  <=    (tmr_registers(0)(109) and tmr_registers(1)(109)) or                                                             
                            (tmr_registers(1)(109) and tmr_registers(2)(109)) or                                                             
                            (tmr_registers(0)(109) and tmr_registers(2)(109));                                                               
                                                                                                                                         
        local_tmr_voter(110)  <=    (tmr_registers(0)(110) and tmr_registers(1)(110)) or                                                             
                            (tmr_registers(1)(110) and tmr_registers(2)(110)) or                                                             
                            (tmr_registers(0)(110) and tmr_registers(2)(110));                                                               
                                                                                                                                         
        local_tmr_voter(111)  <=    (tmr_registers(0)(111) and tmr_registers(1)(111)) or                                                             
                            (tmr_registers(1)(111) and tmr_registers(2)(111)) or                                                             
                            (tmr_registers(0)(111) and tmr_registers(2)(111));                                                               
                                                                                                                                         
        local_tmr_voter(112)  <=    (tmr_registers(0)(112) and tmr_registers(1)(112)) or                                                             
                            (tmr_registers(1)(112) and tmr_registers(2)(112)) or                                                             
                            (tmr_registers(0)(112) and tmr_registers(2)(112));                                                               
                                                                                                                                         
        local_tmr_voter(113)  <=    (tmr_registers(0)(113) and tmr_registers(1)(113)) or                                                             
                            (tmr_registers(1)(113) and tmr_registers(2)(113)) or                                                             
                            (tmr_registers(0)(113) and tmr_registers(2)(113));                                                               
                                                                                                                                         
        local_tmr_voter(114)  <=    (tmr_registers(0)(114) and tmr_registers(1)(114)) or                                                             
                            (tmr_registers(1)(114) and tmr_registers(2)(114)) or                                                             
                            (tmr_registers(0)(114) and tmr_registers(2)(114));                                                               
                                                                                                                                         
        local_tmr_voter(115)  <=    (tmr_registers(0)(115) and tmr_registers(1)(115)) or                                                             
                            (tmr_registers(1)(115) and tmr_registers(2)(115)) or                                                             
                            (tmr_registers(0)(115) and tmr_registers(2)(115));                                                               
                                                                                                                                         
        local_tmr_voter(116)  <=    (tmr_registers(0)(116) and tmr_registers(1)(116)) or                                                             
                            (tmr_registers(1)(116) and tmr_registers(2)(116)) or                                                             
                            (tmr_registers(0)(116) and tmr_registers(2)(116));                                                               
                                                                                                                                         
        local_tmr_voter(117)  <=    (tmr_registers(0)(117) and tmr_registers(1)(117)) or                                                             
                            (tmr_registers(1)(117) and tmr_registers(2)(117)) or                                                             
                            (tmr_registers(0)(117) and tmr_registers(2)(117));                                                               
                                                                                                                                         
        local_tmr_voter(118)  <=    (tmr_registers(0)(118) and tmr_registers(1)(118)) or                                                             
                            (tmr_registers(1)(118) and tmr_registers(2)(118)) or                                                             
                            (tmr_registers(0)(118) and tmr_registers(2)(118));                                                               
                                                                                                                                         
        local_tmr_voter(119)  <=    (tmr_registers(0)(119) and tmr_registers(1)(119)) or                                                             
                            (tmr_registers(1)(119) and tmr_registers(2)(119)) or                                                             
                            (tmr_registers(0)(119) and tmr_registers(2)(119));                                                               
                                                                                                                                         
        local_tmr_voter(120)  <=    (tmr_registers(0)(120) and tmr_registers(1)(120)) or                                                             
                            (tmr_registers(1)(120) and tmr_registers(2)(120)) or                                                             
                            (tmr_registers(0)(120) and tmr_registers(2)(120));                                                               
                                                                                                                                         
        local_tmr_voter(121)  <=    (tmr_registers(0)(121) and tmr_registers(1)(121)) or                                                             
                            (tmr_registers(1)(121) and tmr_registers(2)(121)) or                                                             
                            (tmr_registers(0)(121) and tmr_registers(2)(121));                                                               
                                                                                                                                         
        local_tmr_voter(122)  <=    (tmr_registers(0)(122) and tmr_registers(1)(122)) or                                                             
                            (tmr_registers(1)(122) and tmr_registers(2)(122)) or                                                             
                            (tmr_registers(0)(122) and tmr_registers(2)(122));                                                               
                                                                                                                                         
        local_tmr_voter(123)  <=    (tmr_registers(0)(123) and tmr_registers(1)(123)) or                                                             
                            (tmr_registers(1)(123) and tmr_registers(2)(123)) or                                                             
                            (tmr_registers(0)(123) and tmr_registers(2)(123));                                                               
                                                                                                                                         
        local_tmr_voter(124)  <=    (tmr_registers(0)(124) and tmr_registers(1)(124)) or                                                             
                            (tmr_registers(1)(124) and tmr_registers(2)(124)) or                                                             
                            (tmr_registers(0)(124) and tmr_registers(2)(124));                                                               
                                                                                                                                         
        local_tmr_voter(125)  <=    (tmr_registers(0)(125) and tmr_registers(1)(125)) or                                                             
                            (tmr_registers(1)(125) and tmr_registers(2)(125)) or                                                             
                            (tmr_registers(0)(125) and tmr_registers(2)(125));                                                               
                                                                                                                                         
        local_tmr_voter(126)  <=    (tmr_registers(0)(126) and tmr_registers(1)(126)) or                                                             
                            (tmr_registers(1)(126) and tmr_registers(2)(126)) or                                                             
                            (tmr_registers(0)(126) and tmr_registers(2)(126));                                                               
                                                                                                                                         
        local_tmr_voter(127)  <=    (tmr_registers(0)(127) and tmr_registers(1)(127)) or                                                             
                            (tmr_registers(1)(127) and tmr_registers(2)(127)) or                                                             
                            (tmr_registers(0)(127) and tmr_registers(2)(127));                                                               
                                                                                                                                         
        local_tmr_voter(128)  <=    (tmr_registers(0)(128) and tmr_registers(1)(128)) or                                                             
                            (tmr_registers(1)(128) and tmr_registers(2)(128)) or                                                             
                            (tmr_registers(0)(128) and tmr_registers(2)(128));                                                               
                                                                                                                                         
        local_tmr_voter(129)  <=    (tmr_registers(0)(129) and tmr_registers(1)(129)) or                                                             
                            (tmr_registers(1)(129) and tmr_registers(2)(129)) or                                                             
                            (tmr_registers(0)(129) and tmr_registers(2)(129));                                                               
                                                                                                                                         
        local_tmr_voter(130)  <=    (tmr_registers(0)(130) and tmr_registers(1)(130)) or                                                             
                            (tmr_registers(1)(130) and tmr_registers(2)(130)) or                                                             
                            (tmr_registers(0)(130) and tmr_registers(2)(130));                                                               
                                                                                                                                         
        local_tmr_voter(131)  <=    (tmr_registers(0)(131) and tmr_registers(1)(131)) or                                                             
                            (tmr_registers(1)(131) and tmr_registers(2)(131)) or                                                             
                            (tmr_registers(0)(131) and tmr_registers(2)(131));                                                               
                                                                                                                                         
        local_tmr_voter(132)  <=    (tmr_registers(0)(132) and tmr_registers(1)(132)) or                                                             
                            (tmr_registers(1)(132) and tmr_registers(2)(132)) or                                                             
                            (tmr_registers(0)(132) and tmr_registers(2)(132));                                                               
                                                                                                                                         
        local_tmr_voter(133)  <=    (tmr_registers(0)(133) and tmr_registers(1)(133)) or                                                             
                            (tmr_registers(1)(133) and tmr_registers(2)(133)) or                                                             
                            (tmr_registers(0)(133) and tmr_registers(2)(133));                                                               
                                                                                                                                         
        local_tmr_voter(134)  <=    (tmr_registers(0)(134) and tmr_registers(1)(134)) or                                                             
                            (tmr_registers(1)(134) and tmr_registers(2)(134)) or                                                             
                            (tmr_registers(0)(134) and tmr_registers(2)(134));                                                               
                                                                                                                                         
        local_tmr_voter(135)  <=    (tmr_registers(0)(135) and tmr_registers(1)(135)) or                                                             
                            (tmr_registers(1)(135) and tmr_registers(2)(135)) or                                                             
                            (tmr_registers(0)(135) and tmr_registers(2)(135));                                                               
                                                                                                                                         
        local_tmr_voter(136)  <=    (tmr_registers(0)(136) and tmr_registers(1)(136)) or                                                             
                            (tmr_registers(1)(136) and tmr_registers(2)(136)) or                                                             
                            (tmr_registers(0)(136) and tmr_registers(2)(136));                                                               
                                                                                                                                         
        local_tmr_voter(137)  <=    (tmr_registers(0)(137) and tmr_registers(1)(137)) or                                                             
                            (tmr_registers(1)(137) and tmr_registers(2)(137)) or                                                             
                            (tmr_registers(0)(137) and tmr_registers(2)(137));                                                               
                                                                                                                                         
        local_tmr_voter(138)  <=    (tmr_registers(0)(138) and tmr_registers(1)(138)) or                                                             
                            (tmr_registers(1)(138) and tmr_registers(2)(138)) or                                                             
                            (tmr_registers(0)(138) and tmr_registers(2)(138));                                                               
                                                                                                                                         
        local_tmr_voter(139)  <=    (tmr_registers(0)(139) and tmr_registers(1)(139)) or                                                             
                            (tmr_registers(1)(139) and tmr_registers(2)(139)) or                                                             
                            (tmr_registers(0)(139) and tmr_registers(2)(139));                                                               
                                                                                                                                         
        local_tmr_voter(140)  <=    (tmr_registers(0)(140) and tmr_registers(1)(140)) or                                                             
                            (tmr_registers(1)(140) and tmr_registers(2)(140)) or                                                             
                            (tmr_registers(0)(140) and tmr_registers(2)(140));                                                               
                                                                                                                                         
        local_tmr_voter(141)  <=    (tmr_registers(0)(141) and tmr_registers(1)(141)) or                                                             
                            (tmr_registers(1)(141) and tmr_registers(2)(141)) or                                                             
                            (tmr_registers(0)(141) and tmr_registers(2)(141));                                                               
                                                                                                                                         
        local_tmr_voter(142)  <=    (tmr_registers(0)(142) and tmr_registers(1)(142)) or                                                             
                            (tmr_registers(1)(142) and tmr_registers(2)(142)) or                                                             
                            (tmr_registers(0)(142) and tmr_registers(2)(142));                                                               
                                                                                                                                         
        local_tmr_voter(143)  <=    (tmr_registers(0)(143) and tmr_registers(1)(143)) or                                                             
                            (tmr_registers(1)(143) and tmr_registers(2)(143)) or                                                             
                            (tmr_registers(0)(143) and tmr_registers(2)(143));                                                               
                                                                                                                                         
        local_tmr_voter(144)  <=    (tmr_registers(0)(144) and tmr_registers(1)(144)) or                                                             
                            (tmr_registers(1)(144) and tmr_registers(2)(144)) or                                                             
                            (tmr_registers(0)(144) and tmr_registers(2)(144));                                                               
                                                                                                                                         
        local_tmr_voter(145)  <=    (tmr_registers(0)(145) and tmr_registers(1)(145)) or                                                             
                            (tmr_registers(1)(145) and tmr_registers(2)(145)) or                                                             
                            (tmr_registers(0)(145) and tmr_registers(2)(145));                                                               
                                                                                                                                         
        local_tmr_voter(146)  <=    (tmr_registers(0)(146) and tmr_registers(1)(146)) or                                                             
                            (tmr_registers(1)(146) and tmr_registers(2)(146)) or                                                             
                            (tmr_registers(0)(146) and tmr_registers(2)(146));                                                               
                                                                                                                                         
        local_tmr_voter(147)  <=    (tmr_registers(0)(147) and tmr_registers(1)(147)) or                                                             
                            (tmr_registers(1)(147) and tmr_registers(2)(147)) or                                                             
                            (tmr_registers(0)(147) and tmr_registers(2)(147));                                                               
                                                                                                                                         
        local_tmr_voter(148)  <=    (tmr_registers(0)(148) and tmr_registers(1)(148)) or                                                             
                            (tmr_registers(1)(148) and tmr_registers(2)(148)) or                                                             
                            (tmr_registers(0)(148) and tmr_registers(2)(148));                                                               
                                                                                                                                         
        local_tmr_voter(149)  <=    (tmr_registers(0)(149) and tmr_registers(1)(149)) or                                                             
                            (tmr_registers(1)(149) and tmr_registers(2)(149)) or                                                             
                            (tmr_registers(0)(149) and tmr_registers(2)(149));                                                               
                                                                                                                                         
        local_tmr_voter(150)  <=    (tmr_registers(0)(150) and tmr_registers(1)(150)) or                                                             
                            (tmr_registers(1)(150) and tmr_registers(2)(150)) or                                                             
                            (tmr_registers(0)(150) and tmr_registers(2)(150));                                                               
                                                                                                                                         
        local_tmr_voter(151)  <=    (tmr_registers(0)(151) and tmr_registers(1)(151)) or                                                             
                            (tmr_registers(1)(151) and tmr_registers(2)(151)) or                                                             
                            (tmr_registers(0)(151) and tmr_registers(2)(151));                                                               
                                                                                                                                         
        local_tmr_voter(152)  <=    (tmr_registers(0)(152) and tmr_registers(1)(152)) or                                                             
                            (tmr_registers(1)(152) and tmr_registers(2)(152)) or                                                             
                            (tmr_registers(0)(152) and tmr_registers(2)(152));                                                               
                                                                                                                                         
        local_tmr_voter(153)  <=    (tmr_registers(0)(153) and tmr_registers(1)(153)) or                                                             
                            (tmr_registers(1)(153) and tmr_registers(2)(153)) or                                                             
                            (tmr_registers(0)(153) and tmr_registers(2)(153));                                                               
                                                                                                                                         
        local_tmr_voter(154)  <=    (tmr_registers(0)(154) and tmr_registers(1)(154)) or                                                             
                            (tmr_registers(1)(154) and tmr_registers(2)(154)) or                                                             
                            (tmr_registers(0)(154) and tmr_registers(2)(154));                                                               
                                                                                                                                         
        local_tmr_voter(155)  <=    (tmr_registers(0)(155) and tmr_registers(1)(155)) or                                                             
                            (tmr_registers(1)(155) and tmr_registers(2)(155)) or                                                             
                            (tmr_registers(0)(155) and tmr_registers(2)(155));                                                               
                                                                                                                                         
        local_tmr_voter(156)  <=    (tmr_registers(0)(156) and tmr_registers(1)(156)) or                                                             
                            (tmr_registers(1)(156) and tmr_registers(2)(156)) or                                                             
                            (tmr_registers(0)(156) and tmr_registers(2)(156));                                                               
                                                                                                                                         
        local_tmr_voter(157)  <=    (tmr_registers(0)(157) and tmr_registers(1)(157)) or                                                             
                            (tmr_registers(1)(157) and tmr_registers(2)(157)) or                                                             
                            (tmr_registers(0)(157) and tmr_registers(2)(157));                                                               
                                                                                                                                         
        local_tmr_voter(158)  <=    (tmr_registers(0)(158) and tmr_registers(1)(158)) or                                                             
                            (tmr_registers(1)(158) and tmr_registers(2)(158)) or                                                             
                            (tmr_registers(0)(158) and tmr_registers(2)(158));                                                               
                                                                                                                                         
        local_tmr_voter(159)  <=    (tmr_registers(0)(159) and tmr_registers(1)(159)) or                                                             
                            (tmr_registers(1)(159) and tmr_registers(2)(159)) or                                                             
                            (tmr_registers(0)(159) and tmr_registers(2)(159));                                                               
                                                                                                                                         
        local_tmr_voter(160)  <=    (tmr_registers(0)(160) and tmr_registers(1)(160)) or                                                             
                            (tmr_registers(1)(160) and tmr_registers(2)(160)) or                                                             
                            (tmr_registers(0)(160) and tmr_registers(2)(160));                                                               
                                                                                                                                         
        local_tmr_voter(161)  <=    (tmr_registers(0)(161) and tmr_registers(1)(161)) or                                                             
                            (tmr_registers(1)(161) and tmr_registers(2)(161)) or                                                             
                            (tmr_registers(0)(161) and tmr_registers(2)(161));                                                               
                                                                                                                                         
        local_tmr_voter(162)  <=    (tmr_registers(0)(162) and tmr_registers(1)(162)) or                                                             
                            (tmr_registers(1)(162) and tmr_registers(2)(162)) or                                                             
                            (tmr_registers(0)(162) and tmr_registers(2)(162));                                                               
                                                                                                                                         
        local_tmr_voter(163)  <=    (tmr_registers(0)(163) and tmr_registers(1)(163)) or                                                             
                            (tmr_registers(1)(163) and tmr_registers(2)(163)) or                                                             
                            (tmr_registers(0)(163) and tmr_registers(2)(163));                                                               
                                                                                                                                         
        local_tmr_voter(164)  <=    (tmr_registers(0)(164) and tmr_registers(1)(164)) or                                                             
                            (tmr_registers(1)(164) and tmr_registers(2)(164)) or                                                             
                            (tmr_registers(0)(164) and tmr_registers(2)(164));                                                               
                                                                                                                                         
        local_tmr_voter(165)  <=    (tmr_registers(0)(165) and tmr_registers(1)(165)) or                                                             
                            (tmr_registers(1)(165) and tmr_registers(2)(165)) or                                                             
                            (tmr_registers(0)(165) and tmr_registers(2)(165));                                                               
                                                                                                                                         
        local_tmr_voter(166)  <=    (tmr_registers(0)(166) and tmr_registers(1)(166)) or                                                             
                            (tmr_registers(1)(166) and tmr_registers(2)(166)) or                                                             
                            (tmr_registers(0)(166) and tmr_registers(2)(166));                                                               
                                                                                                                                         
        local_tmr_voter(167)  <=    (tmr_registers(0)(167) and tmr_registers(1)(167)) or                                                             
                            (tmr_registers(1)(167) and tmr_registers(2)(167)) or                                                             
                            (tmr_registers(0)(167) and tmr_registers(2)(167));                                                               
                                                                                                                                         
        local_tmr_voter(168)  <=    (tmr_registers(0)(168) and tmr_registers(1)(168)) or                                                             
                            (tmr_registers(1)(168) and tmr_registers(2)(168)) or                                                             
                            (tmr_registers(0)(168) and tmr_registers(2)(168));                                                               
                                                                                                                                         
        local_tmr_voter(169)  <=    (tmr_registers(0)(169) and tmr_registers(1)(169)) or                                                             
                            (tmr_registers(1)(169) and tmr_registers(2)(169)) or                                                             
                            (tmr_registers(0)(169) and tmr_registers(2)(169));                                                               
                                                                                                                                         
        local_tmr_voter(170)  <=    (tmr_registers(0)(170) and tmr_registers(1)(170)) or                                                             
                            (tmr_registers(1)(170) and tmr_registers(2)(170)) or                                                             
                            (tmr_registers(0)(170) and tmr_registers(2)(170));                                                               
                                                                                                                                         
        local_tmr_voter(171)  <=    (tmr_registers(0)(171) and tmr_registers(1)(171)) or                                                             
                            (tmr_registers(1)(171) and tmr_registers(2)(171)) or                                                             
                            (tmr_registers(0)(171) and tmr_registers(2)(171));                                                               
                                                                                                                                         
        local_tmr_voter(172)  <=    (tmr_registers(0)(172) and tmr_registers(1)(172)) or                                                             
                            (tmr_registers(1)(172) and tmr_registers(2)(172)) or                                                             
                            (tmr_registers(0)(172) and tmr_registers(2)(172));                                                               
                                                                                                                                         
        local_tmr_voter(173)  <=    (tmr_registers(0)(173) and tmr_registers(1)(173)) or                                                             
                            (tmr_registers(1)(173) and tmr_registers(2)(173)) or                                                             
                            (tmr_registers(0)(173) and tmr_registers(2)(173));                                                               
                                                                                                                                         
        local_tmr_voter(174)  <=    (tmr_registers(0)(174) and tmr_registers(1)(174)) or                                                             
                            (tmr_registers(1)(174) and tmr_registers(2)(174)) or                                                             
                            (tmr_registers(0)(174) and tmr_registers(2)(174));                                                               
                                                                                                                                         
        local_tmr_voter(175)  <=    (tmr_registers(0)(175) and tmr_registers(1)(175)) or                                                             
                            (tmr_registers(1)(175) and tmr_registers(2)(175)) or                                                             
                            (tmr_registers(0)(175) and tmr_registers(2)(175));                                                               
                                                                                                                                         
        local_tmr_voter(176)  <=    (tmr_registers(0)(176) and tmr_registers(1)(176)) or                                                             
                            (tmr_registers(1)(176) and tmr_registers(2)(176)) or                                                             
                            (tmr_registers(0)(176) and tmr_registers(2)(176));                                                               
                                                                                                                                         
        local_tmr_voter(177)  <=    (tmr_registers(0)(177) and tmr_registers(1)(177)) or                                                             
                            (tmr_registers(1)(177) and tmr_registers(2)(177)) or                                                             
                            (tmr_registers(0)(177) and tmr_registers(2)(177));                                                               
                                                                                                                                         
        local_tmr_voter(178)  <=    (tmr_registers(0)(178) and tmr_registers(1)(178)) or                                                             
                            (tmr_registers(1)(178) and tmr_registers(2)(178)) or                                                             
                            (tmr_registers(0)(178) and tmr_registers(2)(178));                                                               
                                                                                                                                         
        local_tmr_voter(179)  <=    (tmr_registers(0)(179) and tmr_registers(1)(179)) or                                                             
                            (tmr_registers(1)(179) and tmr_registers(2)(179)) or                                                             
                            (tmr_registers(0)(179) and tmr_registers(2)(179));                                                               
                                                                                                                                         
        local_tmr_voter(180)  <=    (tmr_registers(0)(180) and tmr_registers(1)(180)) or                                                             
                            (tmr_registers(1)(180) and tmr_registers(2)(180)) or                                                             
                            (tmr_registers(0)(180) and tmr_registers(2)(180));                                                               
                                                                                                                                         
        local_tmr_voter(181)  <=    (tmr_registers(0)(181) and tmr_registers(1)(181)) or                                                             
                            (tmr_registers(1)(181) and tmr_registers(2)(181)) or                                                             
                            (tmr_registers(0)(181) and tmr_registers(2)(181));                                                               
                                                                                                                                         
        local_tmr_voter(182)  <=    (tmr_registers(0)(182) and tmr_registers(1)(182)) or                                                             
                            (tmr_registers(1)(182) and tmr_registers(2)(182)) or                                                             
                            (tmr_registers(0)(182) and tmr_registers(2)(182));                                                               
                                                                                                                                         
        local_tmr_voter(183)  <=    (tmr_registers(0)(183) and tmr_registers(1)(183)) or                                                             
                            (tmr_registers(1)(183) and tmr_registers(2)(183)) or                                                             
                            (tmr_registers(0)(183) and tmr_registers(2)(183));                                                               
                                                                                                                                         
        local_tmr_voter(184)  <=    (tmr_registers(0)(184) and tmr_registers(1)(184)) or                                                             
                            (tmr_registers(1)(184) and tmr_registers(2)(184)) or                                                             
                            (tmr_registers(0)(184) and tmr_registers(2)(184));                                                               
                                                                                                                                         
        local_tmr_voter(185)  <=    (tmr_registers(0)(185) and tmr_registers(1)(185)) or                                                             
                            (tmr_registers(1)(185) and tmr_registers(2)(185)) or                                                             
                            (tmr_registers(0)(185) and tmr_registers(2)(185));                                                               
                                                                                                                                         
        local_tmr_voter(186)  <=    (tmr_registers(0)(186) and tmr_registers(1)(186)) or                                                             
                            (tmr_registers(1)(186) and tmr_registers(2)(186)) or                                                             
                            (tmr_registers(0)(186) and tmr_registers(2)(186));                                                               
                                                                                                                                         
        local_tmr_voter(187)  <=    (tmr_registers(0)(187) and tmr_registers(1)(187)) or                                                             
                            (tmr_registers(1)(187) and tmr_registers(2)(187)) or                                                             
                            (tmr_registers(0)(187) and tmr_registers(2)(187));                                                               
                                                                                                                                         
        local_tmr_voter(188)  <=    (tmr_registers(0)(188) and tmr_registers(1)(188)) or                                                             
                            (tmr_registers(1)(188) and tmr_registers(2)(188)) or                                                             
                            (tmr_registers(0)(188) and tmr_registers(2)(188));                                                               
                                                                                                                                         
        local_tmr_voter(189)  <=    (tmr_registers(0)(189) and tmr_registers(1)(189)) or                                                             
                            (tmr_registers(1)(189) and tmr_registers(2)(189)) or                                                             
                            (tmr_registers(0)(189) and tmr_registers(2)(189));                                                               
                                                                                                                                         
        local_tmr_voter(190)  <=    (tmr_registers(0)(190) and tmr_registers(1)(190)) or                                                             
                            (tmr_registers(1)(190) and tmr_registers(2)(190)) or                                                             
                            (tmr_registers(0)(190) and tmr_registers(2)(190));                                                               
                                                                                                                                         
        local_tmr_voter(191)  <=    (tmr_registers(0)(191) and tmr_registers(1)(191)) or                                                             
                            (tmr_registers(1)(191) and tmr_registers(2)(191)) or                                                             
                            (tmr_registers(0)(191) and tmr_registers(2)(191));                                                               
                                                                                                                                         
        local_tmr_voter(192)  <=    (tmr_registers(0)(192) and tmr_registers(1)(192)) or                                                             
                            (tmr_registers(1)(192) and tmr_registers(2)(192)) or                                                             
                            (tmr_registers(0)(192) and tmr_registers(2)(192));                                                               
                                                                                                                                         
        local_tmr_voter(193)  <=    (tmr_registers(0)(193) and tmr_registers(1)(193)) or                                                             
                            (tmr_registers(1)(193) and tmr_registers(2)(193)) or                                                             
                            (tmr_registers(0)(193) and tmr_registers(2)(193));                                                               
                                                                                                                                         
        local_tmr_voter(194)  <=    (tmr_registers(0)(194) and tmr_registers(1)(194)) or                                                             
                            (tmr_registers(1)(194) and tmr_registers(2)(194)) or                                                             
                            (tmr_registers(0)(194) and tmr_registers(2)(194));                                                               
                                                                                                                                         
        local_tmr_voter(195)  <=    (tmr_registers(0)(195) and tmr_registers(1)(195)) or                                                             
                            (tmr_registers(1)(195) and tmr_registers(2)(195)) or                                                             
                            (tmr_registers(0)(195) and tmr_registers(2)(195));                                                               
                                                                                                                                         
        local_tmr_voter(196)  <=    (tmr_registers(0)(196) and tmr_registers(1)(196)) or                                                             
                            (tmr_registers(1)(196) and tmr_registers(2)(196)) or                                                             
                            (tmr_registers(0)(196) and tmr_registers(2)(196));                                                               
                                                                                                                                         
        local_tmr_voter(197)  <=    (tmr_registers(0)(197) and tmr_registers(1)(197)) or                                                             
                            (tmr_registers(1)(197) and tmr_registers(2)(197)) or                                                             
                            (tmr_registers(0)(197) and tmr_registers(2)(197));                                                               
                                                                                                                                         
        local_tmr_voter(198)  <=    (tmr_registers(0)(198) and tmr_registers(1)(198)) or                                                             
                            (tmr_registers(1)(198) and tmr_registers(2)(198)) or                                                             
                            (tmr_registers(0)(198) and tmr_registers(2)(198));                                                               
                                                                                                                                         
        local_tmr_voter(199)  <=    (tmr_registers(0)(199) and tmr_registers(1)(199)) or                                                             
                            (tmr_registers(1)(199) and tmr_registers(2)(199)) or                                                             
                            (tmr_registers(0)(199) and tmr_registers(2)(199));                                                               
                                                                                                                                         
        local_tmr_voter(200)  <=    (tmr_registers(0)(200) and tmr_registers(1)(200)) or                                                             
                            (tmr_registers(1)(200) and tmr_registers(2)(200)) or                                                             
                            (tmr_registers(0)(200) and tmr_registers(2)(200));                                                               
                                                                                                                                         
        local_tmr_voter(201)  <=    (tmr_registers(0)(201) and tmr_registers(1)(201)) or                                                             
                            (tmr_registers(1)(201) and tmr_registers(2)(201)) or                                                             
                            (tmr_registers(0)(201) and tmr_registers(2)(201));                                                               
                                                                                                                                         
        local_tmr_voter(202)  <=    (tmr_registers(0)(202) and tmr_registers(1)(202)) or                                                             
                            (tmr_registers(1)(202) and tmr_registers(2)(202)) or                                                             
                            (tmr_registers(0)(202) and tmr_registers(2)(202));                                                               
                                                                                                                                         
        local_tmr_voter(203)  <=    (tmr_registers(0)(203) and tmr_registers(1)(203)) or                                                             
                            (tmr_registers(1)(203) and tmr_registers(2)(203)) or                                                             
                            (tmr_registers(0)(203) and tmr_registers(2)(203));                                                               
                                                                                                                                         
        local_tmr_voter(204)  <=    (tmr_registers(0)(204) and tmr_registers(1)(204)) or                                                             
                            (tmr_registers(1)(204) and tmr_registers(2)(204)) or                                                             
                            (tmr_registers(0)(204) and tmr_registers(2)(204));                                                               
                                                                                                                                         
        local_tmr_voter(205)  <=    (tmr_registers(0)(205) and tmr_registers(1)(205)) or                                                             
                            (tmr_registers(1)(205) and tmr_registers(2)(205)) or                                                             
                            (tmr_registers(0)(205) and tmr_registers(2)(205));                                                               
                                                                                                                                         
        local_tmr_voter(206)  <=    (tmr_registers(0)(206) and tmr_registers(1)(206)) or                                                             
                            (tmr_registers(1)(206) and tmr_registers(2)(206)) or                                                             
                            (tmr_registers(0)(206) and tmr_registers(2)(206));                                                               
                                                                                                                                         
        local_tmr_voter(207)  <=    (tmr_registers(0)(207) and tmr_registers(1)(207)) or                                                             
                            (tmr_registers(1)(207) and tmr_registers(2)(207)) or                                                             
                            (tmr_registers(0)(207) and tmr_registers(2)(207));                                                               
                                                                                                                                         
        local_tmr_voter(208)  <=    (tmr_registers(0)(208) and tmr_registers(1)(208)) or                                                             
                            (tmr_registers(1)(208) and tmr_registers(2)(208)) or                                                             
                            (tmr_registers(0)(208) and tmr_registers(2)(208));                                                               
                                                                                                                                         
        local_tmr_voter(209)  <=    (tmr_registers(0)(209) and tmr_registers(1)(209)) or                                                             
                            (tmr_registers(1)(209) and tmr_registers(2)(209)) or                                                             
                            (tmr_registers(0)(209) and tmr_registers(2)(209));                                                               
                                                                                                                                         
        local_tmr_voter(210)  <=    (tmr_registers(0)(210) and tmr_registers(1)(210)) or                                                             
                            (tmr_registers(1)(210) and tmr_registers(2)(210)) or                                                             
                            (tmr_registers(0)(210) and tmr_registers(2)(210));                                                               
                                                                                                                                         
        local_tmr_voter(211)  <=    (tmr_registers(0)(211) and tmr_registers(1)(211)) or                                                             
                            (tmr_registers(1)(211) and tmr_registers(2)(211)) or                                                             
                            (tmr_registers(0)(211) and tmr_registers(2)(211));                                                               
                                                                                                                                         
        local_tmr_voter(212)  <=    (tmr_registers(0)(212) and tmr_registers(1)(212)) or                                                             
                            (tmr_registers(1)(212) and tmr_registers(2)(212)) or                                                             
                            (tmr_registers(0)(212) and tmr_registers(2)(212));                                                               
                                                                                                                                         
        local_tmr_voter(213)  <=    (tmr_registers(0)(213) and tmr_registers(1)(213)) or                                                             
                            (tmr_registers(1)(213) and tmr_registers(2)(213)) or                                                             
                            (tmr_registers(0)(213) and tmr_registers(2)(213));                                                               
                                                                                                                                         
        local_tmr_voter(214)  <=    (tmr_registers(0)(214) and tmr_registers(1)(214)) or                                                             
                            (tmr_registers(1)(214) and tmr_registers(2)(214)) or                                                             
                            (tmr_registers(0)(214) and tmr_registers(2)(214));                                                               
                                                                                                                                         
        local_tmr_voter(215)  <=    (tmr_registers(0)(215) and tmr_registers(1)(215)) or                                                             
                            (tmr_registers(1)(215) and tmr_registers(2)(215)) or                                                             
                            (tmr_registers(0)(215) and tmr_registers(2)(215));                                                               
                                                                                                                                         
        local_tmr_voter(216)  <=    (tmr_registers(0)(216) and tmr_registers(1)(216)) or                                                             
                            (tmr_registers(1)(216) and tmr_registers(2)(216)) or                                                             
                            (tmr_registers(0)(216) and tmr_registers(2)(216));                                                               
                                                                                                                                         
        local_tmr_voter(217)  <=    (tmr_registers(0)(217) and tmr_registers(1)(217)) or                                                             
                            (tmr_registers(1)(217) and tmr_registers(2)(217)) or                                                             
                            (tmr_registers(0)(217) and tmr_registers(2)(217));                                                               
                                                                                                                                         
        local_tmr_voter(218)  <=    (tmr_registers(0)(218) and tmr_registers(1)(218)) or                                                             
                            (tmr_registers(1)(218) and tmr_registers(2)(218)) or                                                             
                            (tmr_registers(0)(218) and tmr_registers(2)(218));                                                               
                                                                                                                                         
        local_tmr_voter(219)  <=    (tmr_registers(0)(219) and tmr_registers(1)(219)) or                                                             
                            (tmr_registers(1)(219) and tmr_registers(2)(219)) or                                                             
                            (tmr_registers(0)(219) and tmr_registers(2)(219));                                                               
                                                                                                                                         
        local_tmr_voter(220)  <=    (tmr_registers(0)(220) and tmr_registers(1)(220)) or                                                             
                            (tmr_registers(1)(220) and tmr_registers(2)(220)) or                                                             
                            (tmr_registers(0)(220) and tmr_registers(2)(220));                                                               
                                                                                                                                         
        local_tmr_voter(221)  <=    (tmr_registers(0)(221) and tmr_registers(1)(221)) or                                                             
                            (tmr_registers(1)(221) and tmr_registers(2)(221)) or                                                             
                            (tmr_registers(0)(221) and tmr_registers(2)(221));                                                               
                                                                                                                                         
        local_tmr_voter(222)  <=    (tmr_registers(0)(222) and tmr_registers(1)(222)) or                                                             
                            (tmr_registers(1)(222) and tmr_registers(2)(222)) or                                                             
                            (tmr_registers(0)(222) and tmr_registers(2)(222));                                                               
                                                                                                                                         
        local_tmr_voter(223)  <=    (tmr_registers(0)(223) and tmr_registers(1)(223)) or                                                             
                            (tmr_registers(1)(223) and tmr_registers(2)(223)) or                                                             
                            (tmr_registers(0)(223) and tmr_registers(2)(223));                                                               
                                                                                                                                         
        local_tmr_voter(224)  <=    (tmr_registers(0)(224) and tmr_registers(1)(224)) or                                                             
                            (tmr_registers(1)(224) and tmr_registers(2)(224)) or                                                             
                            (tmr_registers(0)(224) and tmr_registers(2)(224));                                                               
                                                                                                                                         
        local_tmr_voter(225)  <=    (tmr_registers(0)(225) and tmr_registers(1)(225)) or                                                             
                            (tmr_registers(1)(225) and tmr_registers(2)(225)) or                                                             
                            (tmr_registers(0)(225) and tmr_registers(2)(225));                                                               
                                                                                                                                         
        local_tmr_voter(226)  <=    (tmr_registers(0)(226) and tmr_registers(1)(226)) or                                                             
                            (tmr_registers(1)(226) and tmr_registers(2)(226)) or                                                             
                            (tmr_registers(0)(226) and tmr_registers(2)(226));                                                               
                                                                                                                                         
        local_tmr_voter(227)  <=    (tmr_registers(0)(227) and tmr_registers(1)(227)) or                                                             
                            (tmr_registers(1)(227) and tmr_registers(2)(227)) or                                                             
                            (tmr_registers(0)(227) and tmr_registers(2)(227));                                                               
                                                                                                                                         
        local_tmr_voter(228)  <=    (tmr_registers(0)(228) and tmr_registers(1)(228)) or                                                             
                            (tmr_registers(1)(228) and tmr_registers(2)(228)) or                                                             
                            (tmr_registers(0)(228) and tmr_registers(2)(228));                                                               
                                                                                                                                         
        local_tmr_voter(229)  <=    (tmr_registers(0)(229) and tmr_registers(1)(229)) or                                                             
                            (tmr_registers(1)(229) and tmr_registers(2)(229)) or                                                             
                            (tmr_registers(0)(229) and tmr_registers(2)(229));                                                               
                                                                                                                                         
        local_tmr_voter(230)  <=    (tmr_registers(0)(230) and tmr_registers(1)(230)) or                                                             
                            (tmr_registers(1)(230) and tmr_registers(2)(230)) or                                                             
                            (tmr_registers(0)(230) and tmr_registers(2)(230));                                                               
                                                                                                                                         
        local_tmr_voter(231)  <=    (tmr_registers(0)(231) and tmr_registers(1)(231)) or                                                             
                            (tmr_registers(1)(231) and tmr_registers(2)(231)) or                                                             
                            (tmr_registers(0)(231) and tmr_registers(2)(231));                                                               
                                                                                                                                         
        local_tmr_voter(232)  <=    (tmr_registers(0)(232) and tmr_registers(1)(232)) or                                                             
                            (tmr_registers(1)(232) and tmr_registers(2)(232)) or                                                             
                            (tmr_registers(0)(232) and tmr_registers(2)(232));                                                               
                                                                                                                                         
        local_tmr_voter(233)  <=    (tmr_registers(0)(233) and tmr_registers(1)(233)) or                                                             
                            (tmr_registers(1)(233) and tmr_registers(2)(233)) or                                                             
                            (tmr_registers(0)(233) and tmr_registers(2)(233));                                                               
                                                                                                                                         
        local_tmr_voter(234)  <=    (tmr_registers(0)(234) and tmr_registers(1)(234)) or                                                             
                            (tmr_registers(1)(234) and tmr_registers(2)(234)) or                                                             
                            (tmr_registers(0)(234) and tmr_registers(2)(234));                                                               
                                                                                                                                         
        local_tmr_voter(235)  <=    (tmr_registers(0)(235) and tmr_registers(1)(235)) or                                                             
                            (tmr_registers(1)(235) and tmr_registers(2)(235)) or                                                             
                            (tmr_registers(0)(235) and tmr_registers(2)(235));                                                               
                                                                                                                                         
        local_tmr_voter(236)  <=    (tmr_registers(0)(236) and tmr_registers(1)(236)) or                                                             
                            (tmr_registers(1)(236) and tmr_registers(2)(236)) or                                                             
                            (tmr_registers(0)(236) and tmr_registers(2)(236));                                                               
                                                                                                                                         
        local_tmr_voter(237)  <=    (tmr_registers(0)(237) and tmr_registers(1)(237)) or                                                             
                            (tmr_registers(1)(237) and tmr_registers(2)(237)) or                                                             
                            (tmr_registers(0)(237) and tmr_registers(2)(237));                                                               
                                                                                                                                         
        local_tmr_voter(238)  <=    (tmr_registers(0)(238) and tmr_registers(1)(238)) or                                                             
                            (tmr_registers(1)(238) and tmr_registers(2)(238)) or                                                             
                            (tmr_registers(0)(238) and tmr_registers(2)(238));                                                               
                                                                                                                                         
        local_tmr_voter(239)  <=    (tmr_registers(0)(239) and tmr_registers(1)(239)) or                                                             
                            (tmr_registers(1)(239) and tmr_registers(2)(239)) or                                                             
                            (tmr_registers(0)(239) and tmr_registers(2)(239));                                                               
                                                                                                                                         
        local_tmr_voter(240)  <=    (tmr_registers(0)(240) and tmr_registers(1)(240)) or                                                             
                            (tmr_registers(1)(240) and tmr_registers(2)(240)) or                                                             
                            (tmr_registers(0)(240) and tmr_registers(2)(240));                                                               
                                                                                                                                         
        local_tmr_voter(241)  <=    (tmr_registers(0)(241) and tmr_registers(1)(241)) or                                                             
                            (tmr_registers(1)(241) and tmr_registers(2)(241)) or                                                             
                            (tmr_registers(0)(241) and tmr_registers(2)(241));                                                               
                                                                                                                                         
        local_tmr_voter(242)  <=    (tmr_registers(0)(242) and tmr_registers(1)(242)) or                                                             
                            (tmr_registers(1)(242) and tmr_registers(2)(242)) or                                                             
                            (tmr_registers(0)(242) and tmr_registers(2)(242));                                                               
                                                                                                                                         
        local_tmr_voter(243)  <=    (tmr_registers(0)(243) and tmr_registers(1)(243)) or                                                             
                            (tmr_registers(1)(243) and tmr_registers(2)(243)) or                                                             
                            (tmr_registers(0)(243) and tmr_registers(2)(243));                                                               
                                                                                                                                         
        local_tmr_voter(244)  <=    (tmr_registers(0)(244) and tmr_registers(1)(244)) or                                                             
                            (tmr_registers(1)(244) and tmr_registers(2)(244)) or                                                             
                            (tmr_registers(0)(244) and tmr_registers(2)(244));                                                               
                                                                                                                                         
        local_tmr_voter(245)  <=    (tmr_registers(0)(245) and tmr_registers(1)(245)) or                                                             
                            (tmr_registers(1)(245) and tmr_registers(2)(245)) or                                                             
                            (tmr_registers(0)(245) and tmr_registers(2)(245));                                                               
                                                                                                                                         
        local_tmr_voter(246)  <=    (tmr_registers(0)(246) and tmr_registers(1)(246)) or                                                             
                            (tmr_registers(1)(246) and tmr_registers(2)(246)) or                                                             
                            (tmr_registers(0)(246) and tmr_registers(2)(246));                                                               
                                                                                                                                         
        local_tmr_voter(247)  <=    (tmr_registers(0)(247) and tmr_registers(1)(247)) or                                                             
                            (tmr_registers(1)(247) and tmr_registers(2)(247)) or                                                             
                            (tmr_registers(0)(247) and tmr_registers(2)(247));                                                               
                                                                                                                                         
        local_tmr_voter(248)  <=    (tmr_registers(0)(248) and tmr_registers(1)(248)) or                                                             
                            (tmr_registers(1)(248) and tmr_registers(2)(248)) or                                                             
                            (tmr_registers(0)(248) and tmr_registers(2)(248));                                                               
                                                                                                                                         
        local_tmr_voter(249)  <=    (tmr_registers(0)(249) and tmr_registers(1)(249)) or                                                             
                            (tmr_registers(1)(249) and tmr_registers(2)(249)) or                                                             
                            (tmr_registers(0)(249) and tmr_registers(2)(249));                                                               
                                                                                                                                         
        local_tmr_voter(250)  <=    (tmr_registers(0)(250) and tmr_registers(1)(250)) or                                                             
                            (tmr_registers(1)(250) and tmr_registers(2)(250)) or                                                             
                            (tmr_registers(0)(250) and tmr_registers(2)(250));                                                               
                                                                                                                                         
        local_tmr_voter(251)  <=    (tmr_registers(0)(251) and tmr_registers(1)(251)) or                                                             
                            (tmr_registers(1)(251) and tmr_registers(2)(251)) or                                                             
                            (tmr_registers(0)(251) and tmr_registers(2)(251));                                                               
                                                                                                                                         
        local_tmr_voter(252)  <=    (tmr_registers(0)(252) and tmr_registers(1)(252)) or                                                             
                            (tmr_registers(1)(252) and tmr_registers(2)(252)) or                                                             
                            (tmr_registers(0)(252) and tmr_registers(2)(252));                                                               
                                                                                                                                         
        local_tmr_voter(253)  <=    (tmr_registers(0)(253) and tmr_registers(1)(253)) or                                                             
                            (tmr_registers(1)(253) and tmr_registers(2)(253)) or                                                             
                            (tmr_registers(0)(253) and tmr_registers(2)(253));                                                               
                                                                                                                                         
        local_tmr_voter(254)  <=    (tmr_registers(0)(254) and tmr_registers(1)(254)) or                                                             
                            (tmr_registers(1)(254) and tmr_registers(2)(254)) or                                                             
                            (tmr_registers(0)(254) and tmr_registers(2)(254));                                                               
                                                                                                                                         
        local_tmr_voter(255)  <=    (tmr_registers(0)(255) and tmr_registers(1)(255)) or                                                             
                            (tmr_registers(1)(255) and tmr_registers(2)(255)) or                                                             
                            (tmr_registers(0)(255) and tmr_registers(2)(255));                                                               
                                                                                                                                         
        local_tmr_voter(256)  <=    (tmr_registers(0)(256) and tmr_registers(1)(256)) or                                                             
                            (tmr_registers(1)(256) and tmr_registers(2)(256)) or                                                             
                            (tmr_registers(0)(256) and tmr_registers(2)(256));                                                               
                                                                                                                                         
        local_tmr_voter(257)  <=    (tmr_registers(0)(257) and tmr_registers(1)(257)) or                                                             
                            (tmr_registers(1)(257) and tmr_registers(2)(257)) or                                                             
                            (tmr_registers(0)(257) and tmr_registers(2)(257));                                                               
                                                                                                                                         
        local_tmr_voter(258)  <=    (tmr_registers(0)(258) and tmr_registers(1)(258)) or                                                             
                            (tmr_registers(1)(258) and tmr_registers(2)(258)) or                                                             
                            (tmr_registers(0)(258) and tmr_registers(2)(258));                                                               
                                                                                                                                         
        local_tmr_voter(259)  <=    (tmr_registers(0)(259) and tmr_registers(1)(259)) or                                                             
                            (tmr_registers(1)(259) and tmr_registers(2)(259)) or                                                             
                            (tmr_registers(0)(259) and tmr_registers(2)(259));                                                               
                                                                                                                                         
        local_tmr_voter(260)  <=    (tmr_registers(0)(260) and tmr_registers(1)(260)) or                                                             
                            (tmr_registers(1)(260) and tmr_registers(2)(260)) or                                                             
                            (tmr_registers(0)(260) and tmr_registers(2)(260));                                                               
                                                                                                                                         
        local_tmr_voter(261)  <=    (tmr_registers(0)(261) and tmr_registers(1)(261)) or                                                             
                            (tmr_registers(1)(261) and tmr_registers(2)(261)) or                                                             
                            (tmr_registers(0)(261) and tmr_registers(2)(261));                                                               
                                                                                                                                         
        local_tmr_voter(262)  <=    (tmr_registers(0)(262) and tmr_registers(1)(262)) or                                                             
                            (tmr_registers(1)(262) and tmr_registers(2)(262)) or                                                             
                            (tmr_registers(0)(262) and tmr_registers(2)(262));                                                               
                                                                                                                                         
        local_tmr_voter(263)  <=    (tmr_registers(0)(263) and tmr_registers(1)(263)) or                                                             
                            (tmr_registers(1)(263) and tmr_registers(2)(263)) or                                                             
                            (tmr_registers(0)(263) and tmr_registers(2)(263));                                                               
                                                                                                                                         
        local_tmr_voter(264)  <=    (tmr_registers(0)(264) and tmr_registers(1)(264)) or                                                             
                            (tmr_registers(1)(264) and tmr_registers(2)(264)) or                                                             
                            (tmr_registers(0)(264) and tmr_registers(2)(264));                                                               
                                                                                                                                         
        local_tmr_voter(265)  <=    (tmr_registers(0)(265) and tmr_registers(1)(265)) or                                                             
                            (tmr_registers(1)(265) and tmr_registers(2)(265)) or                                                             
                            (tmr_registers(0)(265) and tmr_registers(2)(265));                                                               
                                                                                                                                         
        local_tmr_voter(266)  <=    (tmr_registers(0)(266) and tmr_registers(1)(266)) or                                                             
                            (tmr_registers(1)(266) and tmr_registers(2)(266)) or                                                             
                            (tmr_registers(0)(266) and tmr_registers(2)(266));                                                               
                                                                                                                                         
        local_tmr_voter(267)  <=    (tmr_registers(0)(267) and tmr_registers(1)(267)) or                                                             
                            (tmr_registers(1)(267) and tmr_registers(2)(267)) or                                                             
                            (tmr_registers(0)(267) and tmr_registers(2)(267));                                                               
                                                                                                                                         
        local_tmr_voter(268)  <=    (tmr_registers(0)(268) and tmr_registers(1)(268)) or                                                             
                            (tmr_registers(1)(268) and tmr_registers(2)(268)) or                                                             
                            (tmr_registers(0)(268) and tmr_registers(2)(268));                                                               
                                                                                                                                         
        local_tmr_voter(269)  <=    (tmr_registers(0)(269) and tmr_registers(1)(269)) or                                                             
                            (tmr_registers(1)(269) and tmr_registers(2)(269)) or                                                             
                            (tmr_registers(0)(269) and tmr_registers(2)(269));                                                               
                                                                                                                                         
        local_tmr_voter(270)  <=    (tmr_registers(0)(270) and tmr_registers(1)(270)) or                                                             
                            (tmr_registers(1)(270) and tmr_registers(2)(270)) or                                                             
                            (tmr_registers(0)(270) and tmr_registers(2)(270));                                                               
                                                                                                                                         
        local_tmr_voter(271)  <=    (tmr_registers(0)(271) and tmr_registers(1)(271)) or                                                             
                            (tmr_registers(1)(271) and tmr_registers(2)(271)) or                                                             
                            (tmr_registers(0)(271) and tmr_registers(2)(271));                                                               
                                                                                                                                         
        local_tmr_voter(272)  <=    (tmr_registers(0)(272) and tmr_registers(1)(272)) or                                                             
                            (tmr_registers(1)(272) and tmr_registers(2)(272)) or                                                             
                            (tmr_registers(0)(272) and tmr_registers(2)(272));                                                               
                                                                                                                                         
        local_tmr_voter(273)  <=    (tmr_registers(0)(273) and tmr_registers(1)(273)) or                                                             
                            (tmr_registers(1)(273) and tmr_registers(2)(273)) or                                                             
                            (tmr_registers(0)(273) and tmr_registers(2)(273));                                                               
                                                                                                                                         
        local_tmr_voter(274)  <=    (tmr_registers(0)(274) and tmr_registers(1)(274)) or                                                             
                            (tmr_registers(1)(274) and tmr_registers(2)(274)) or                                                             
                            (tmr_registers(0)(274) and tmr_registers(2)(274));                                                               
                                                                                                                                         
        local_tmr_voter(275)  <=    (tmr_registers(0)(275) and tmr_registers(1)(275)) or                                                             
                            (tmr_registers(1)(275) and tmr_registers(2)(275)) or                                                             
                            (tmr_registers(0)(275) and tmr_registers(2)(275));                                                               
                                                                                                                                         
        local_tmr_voter(276)  <=    (tmr_registers(0)(276) and tmr_registers(1)(276)) or                                                             
                            (tmr_registers(1)(276) and tmr_registers(2)(276)) or                                                             
                            (tmr_registers(0)(276) and tmr_registers(2)(276));                                                               
                                                                                                                                         
        local_tmr_voter(277)  <=    (tmr_registers(0)(277) and tmr_registers(1)(277)) or                                                             
                            (tmr_registers(1)(277) and tmr_registers(2)(277)) or                                                             
                            (tmr_registers(0)(277) and tmr_registers(2)(277));                                                               
                                                                                                                                         
        local_tmr_voter(278)  <=    (tmr_registers(0)(278) and tmr_registers(1)(278)) or                                                             
                            (tmr_registers(1)(278) and tmr_registers(2)(278)) or                                                             
                            (tmr_registers(0)(278) and tmr_registers(2)(278));                                                               
                                                                                                                                         
        local_tmr_voter(279)  <=    (tmr_registers(0)(279) and tmr_registers(1)(279)) or                                                             
                            (tmr_registers(1)(279) and tmr_registers(2)(279)) or                                                             
                            (tmr_registers(0)(279) and tmr_registers(2)(279));                                                               
                                                                                                                                         
        local_tmr_voter(280)  <=    (tmr_registers(0)(280) and tmr_registers(1)(280)) or                                                             
                            (tmr_registers(1)(280) and tmr_registers(2)(280)) or                                                             
                            (tmr_registers(0)(280) and tmr_registers(2)(280));                                                               
                                                                                                                                         
        local_tmr_voter(281)  <=    (tmr_registers(0)(281) and tmr_registers(1)(281)) or                                                             
                            (tmr_registers(1)(281) and tmr_registers(2)(281)) or                                                             
                            (tmr_registers(0)(281) and tmr_registers(2)(281));                                                               
                                                                                                                                         
        local_tmr_voter(282)  <=    (tmr_registers(0)(282) and tmr_registers(1)(282)) or                                                             
                            (tmr_registers(1)(282) and tmr_registers(2)(282)) or                                                             
                            (tmr_registers(0)(282) and tmr_registers(2)(282));                                                               
                                                                                                                                         
        local_tmr_voter(283)  <=    (tmr_registers(0)(283) and tmr_registers(1)(283)) or                                                             
                            (tmr_registers(1)(283) and tmr_registers(2)(283)) or                                                             
                            (tmr_registers(0)(283) and tmr_registers(2)(283));                                                               
                                                                                                                                         
        local_tmr_voter(284)  <=    (tmr_registers(0)(284) and tmr_registers(1)(284)) or                                                             
                            (tmr_registers(1)(284) and tmr_registers(2)(284)) or                                                             
                            (tmr_registers(0)(284) and tmr_registers(2)(284));                                                               
                                                                                                                                         
        local_tmr_voter(285)  <=    (tmr_registers(0)(285) and tmr_registers(1)(285)) or                                                             
                            (tmr_registers(1)(285) and tmr_registers(2)(285)) or                                                             
                            (tmr_registers(0)(285) and tmr_registers(2)(285));                                                               
                                                                                                                                         
        local_tmr_voter(286)  <=    (tmr_registers(0)(286) and tmr_registers(1)(286)) or                                                             
                            (tmr_registers(1)(286) and tmr_registers(2)(286)) or                                                             
                            (tmr_registers(0)(286) and tmr_registers(2)(286));                                                               
                                                                                                                                         
        local_tmr_voter(287)  <=    (tmr_registers(0)(287) and tmr_registers(1)(287)) or                                                             
                            (tmr_registers(1)(287) and tmr_registers(2)(287)) or                                                             
                            (tmr_registers(0)(287) and tmr_registers(2)(287));                                                               
                                                                                                                                         
        local_tmr_voter(288)  <=    (tmr_registers(0)(288) and tmr_registers(1)(288)) or                                                             
                            (tmr_registers(1)(288) and tmr_registers(2)(288)) or                                                             
                            (tmr_registers(0)(288) and tmr_registers(2)(288));                                                               
                                                                                                                                         
        local_tmr_voter(289)  <=    (tmr_registers(0)(289) and tmr_registers(1)(289)) or                                                             
                            (tmr_registers(1)(289) and tmr_registers(2)(289)) or                                                             
                            (tmr_registers(0)(289) and tmr_registers(2)(289));                                                               
                                                                                                                                         
        local_tmr_voter(290)  <=    (tmr_registers(0)(290) and tmr_registers(1)(290)) or                                                             
                            (tmr_registers(1)(290) and tmr_registers(2)(290)) or                                                             
                            (tmr_registers(0)(290) and tmr_registers(2)(290));                                                               
                                                                                                                                         
        local_tmr_voter(291)  <=    (tmr_registers(0)(291) and tmr_registers(1)(291)) or                                                             
                            (tmr_registers(1)(291) and tmr_registers(2)(291)) or                                                             
                            (tmr_registers(0)(291) and tmr_registers(2)(291));                                                               
                                                                                                                                         
        local_tmr_voter(292)  <=    (tmr_registers(0)(292) and tmr_registers(1)(292)) or                                                             
                            (tmr_registers(1)(292) and tmr_registers(2)(292)) or                                                             
                            (tmr_registers(0)(292) and tmr_registers(2)(292));                                                               
                                                                                                                                         
        local_tmr_voter(293)  <=    (tmr_registers(0)(293) and tmr_registers(1)(293)) or                                                             
                            (tmr_registers(1)(293) and tmr_registers(2)(293)) or                                                             
                            (tmr_registers(0)(293) and tmr_registers(2)(293));                                                               
                                                                                                                                         
        local_tmr_voter(294)  <=    (tmr_registers(0)(294) and tmr_registers(1)(294)) or                                                             
                            (tmr_registers(1)(294) and tmr_registers(2)(294)) or                                                             
                            (tmr_registers(0)(294) and tmr_registers(2)(294));                                                               
                                                                                                                                         
        local_tmr_voter(295)  <=    (tmr_registers(0)(295) and tmr_registers(1)(295)) or                                                             
                            (tmr_registers(1)(295) and tmr_registers(2)(295)) or                                                             
                            (tmr_registers(0)(295) and tmr_registers(2)(295));                                                               
                                                                                                                                         
        local_tmr_voter(296)  <=    (tmr_registers(0)(296) and tmr_registers(1)(296)) or                                                             
                            (tmr_registers(1)(296) and tmr_registers(2)(296)) or                                                             
                            (tmr_registers(0)(296) and tmr_registers(2)(296));                                                               
                                                                                                                                         
        local_tmr_voter(297)  <=    (tmr_registers(0)(297) and tmr_registers(1)(297)) or                                                             
                            (tmr_registers(1)(297) and tmr_registers(2)(297)) or                                                             
                            (tmr_registers(0)(297) and tmr_registers(2)(297));                                                               
                                                                                                                                         
        local_tmr_voter(298)  <=    (tmr_registers(0)(298) and tmr_registers(1)(298)) or                                                             
                            (tmr_registers(1)(298) and tmr_registers(2)(298)) or                                                             
                            (tmr_registers(0)(298) and tmr_registers(2)(298));                                                               
                                                                                                                                         
        local_tmr_voter(299)  <=    (tmr_registers(0)(299) and tmr_registers(1)(299)) or                                                             
                            (tmr_registers(1)(299) and tmr_registers(2)(299)) or                                                             
                            (tmr_registers(0)(299) and tmr_registers(2)(299));                                                               
                                                                                                                                         
        local_tmr_voter(300)  <=    (tmr_registers(0)(300) and tmr_registers(1)(300)) or                                                             
                            (tmr_registers(1)(300) and tmr_registers(2)(300)) or                                                             
                            (tmr_registers(0)(300) and tmr_registers(2)(300));                                                               
                                                                                                                                         
        local_tmr_voter(301)  <=    (tmr_registers(0)(301) and tmr_registers(1)(301)) or                                                             
                            (tmr_registers(1)(301) and tmr_registers(2)(301)) or                                                             
                            (tmr_registers(0)(301) and tmr_registers(2)(301));                                                               
                                                                                                                                         
        local_tmr_voter(302)  <=    (tmr_registers(0)(302) and tmr_registers(1)(302)) or                                                             
                            (tmr_registers(1)(302) and tmr_registers(2)(302)) or                                                             
                            (tmr_registers(0)(302) and tmr_registers(2)(302));                                                               
                                                                                                                                         
        local_tmr_voter(303)  <=    (tmr_registers(0)(303) and tmr_registers(1)(303)) or                                                             
                            (tmr_registers(1)(303) and tmr_registers(2)(303)) or                                                             
                            (tmr_registers(0)(303) and tmr_registers(2)(303));                                                               
                                                                                                                                         
        local_tmr_voter(304)  <=    (tmr_registers(0)(304) and tmr_registers(1)(304)) or                                                             
                            (tmr_registers(1)(304) and tmr_registers(2)(304)) or                                                             
                            (tmr_registers(0)(304) and tmr_registers(2)(304));                                                               
                                                                                                                                         
        local_tmr_voter(305)  <=    (tmr_registers(0)(305) and tmr_registers(1)(305)) or                                                             
                            (tmr_registers(1)(305) and tmr_registers(2)(305)) or                                                             
                            (tmr_registers(0)(305) and tmr_registers(2)(305));                                                               
                                                                                                                                         
        local_tmr_voter(306)  <=    (tmr_registers(0)(306) and tmr_registers(1)(306)) or                                                             
                            (tmr_registers(1)(306) and tmr_registers(2)(306)) or                                                             
                            (tmr_registers(0)(306) and tmr_registers(2)(306));                                                               
                                                                                                                                         
        local_tmr_voter(307)  <=    (tmr_registers(0)(307) and tmr_registers(1)(307)) or                                                             
                            (tmr_registers(1)(307) and tmr_registers(2)(307)) or                                                             
                            (tmr_registers(0)(307) and tmr_registers(2)(307));                                                               
                                                                                                                                         
        local_tmr_voter(308)  <=    (tmr_registers(0)(308) and tmr_registers(1)(308)) or                                                             
                            (tmr_registers(1)(308) and tmr_registers(2)(308)) or                                                             
                            (tmr_registers(0)(308) and tmr_registers(2)(308));                                                               
                                                                                                                                         
        local_tmr_voter(309)  <=    (tmr_registers(0)(309) and tmr_registers(1)(309)) or                                                             
                            (tmr_registers(1)(309) and tmr_registers(2)(309)) or                                                             
                            (tmr_registers(0)(309) and tmr_registers(2)(309));                                                               
                                                                                                                                         
        local_tmr_voter(310)  <=    (tmr_registers(0)(310) and tmr_registers(1)(310)) or                                                             
                            (tmr_registers(1)(310) and tmr_registers(2)(310)) or                                                             
                            (tmr_registers(0)(310) and tmr_registers(2)(310));                                                               
                                                                                                                                         
        local_tmr_voter(311)  <=    (tmr_registers(0)(311) and tmr_registers(1)(311)) or                                                             
                            (tmr_registers(1)(311) and tmr_registers(2)(311)) or                                                             
                            (tmr_registers(0)(311) and tmr_registers(2)(311));                                                               
                                                                                                                                         
        local_tmr_voter(312)  <=    (tmr_registers(0)(312) and tmr_registers(1)(312)) or                                                             
                            (tmr_registers(1)(312) and tmr_registers(2)(312)) or                                                             
                            (tmr_registers(0)(312) and tmr_registers(2)(312));                                                               
                                                                                                                                         
        local_tmr_voter(313)  <=    (tmr_registers(0)(313) and tmr_registers(1)(313)) or                                                             
                            (tmr_registers(1)(313) and tmr_registers(2)(313)) or                                                             
                            (tmr_registers(0)(313) and tmr_registers(2)(313));                                                               
                                                                                                                                         
        local_tmr_voter(314)  <=    (tmr_registers(0)(314) and tmr_registers(1)(314)) or                                                             
                            (tmr_registers(1)(314) and tmr_registers(2)(314)) or                                                             
                            (tmr_registers(0)(314) and tmr_registers(2)(314));                                                               
                                                                                                                                         
        local_tmr_voter(315)  <=    (tmr_registers(0)(315) and tmr_registers(1)(315)) or                                                             
                            (tmr_registers(1)(315) and tmr_registers(2)(315)) or                                                             
                            (tmr_registers(0)(315) and tmr_registers(2)(315));                                                               
                                                                                                                                         
        local_tmr_voter(316)  <=    (tmr_registers(0)(316) and tmr_registers(1)(316)) or                                                             
                            (tmr_registers(1)(316) and tmr_registers(2)(316)) or                                                             
                            (tmr_registers(0)(316) and tmr_registers(2)(316));                                                               
                                                                                                                                         
        local_tmr_voter(317)  <=    (tmr_registers(0)(317) and tmr_registers(1)(317)) or                                                             
                            (tmr_registers(1)(317) and tmr_registers(2)(317)) or                                                             
                            (tmr_registers(0)(317) and tmr_registers(2)(317));                                                               
                                                                                                                                         
        local_tmr_voter(318)  <=    (tmr_registers(0)(318) and tmr_registers(1)(318)) or                                                             
                            (tmr_registers(1)(318) and tmr_registers(2)(318)) or                                                             
                            (tmr_registers(0)(318) and tmr_registers(2)(318));                                                               
                                                                                                                                         
        local_tmr_voter(319)  <=    (tmr_registers(0)(319) and tmr_registers(1)(319)) or                                                             
                            (tmr_registers(1)(319) and tmr_registers(2)(319)) or                                                             
                            (tmr_registers(0)(319) and tmr_registers(2)(319));                                                               
                                                                                                                                         
        local_tmr_voter(320)  <=    (tmr_registers(0)(320) and tmr_registers(1)(320)) or                                                             
                            (tmr_registers(1)(320) and tmr_registers(2)(320)) or                                                             
                            (tmr_registers(0)(320) and tmr_registers(2)(320));                                                               
                                                                                                                                         
        local_tmr_voter(321)  <=    (tmr_registers(0)(321) and tmr_registers(1)(321)) or                                                             
                            (tmr_registers(1)(321) and tmr_registers(2)(321)) or                                                             
                            (tmr_registers(0)(321) and tmr_registers(2)(321));                                                               
                                                                                                                                         
        local_tmr_voter(322)  <=    (tmr_registers(0)(322) and tmr_registers(1)(322)) or                                                             
                            (tmr_registers(1)(322) and tmr_registers(2)(322)) or                                                             
                            (tmr_registers(0)(322) and tmr_registers(2)(322));                                                               
                                                                                                                                         
        local_tmr_voter(323)  <=    (tmr_registers(0)(323) and tmr_registers(1)(323)) or                                                             
                            (tmr_registers(1)(323) and tmr_registers(2)(323)) or                                                             
                            (tmr_registers(0)(323) and tmr_registers(2)(323));                                                               
                                                                                                                                         
        local_tmr_voter(324)  <=    (tmr_registers(0)(324) and tmr_registers(1)(324)) or                                                             
                            (tmr_registers(1)(324) and tmr_registers(2)(324)) or                                                             
                            (tmr_registers(0)(324) and tmr_registers(2)(324));                                                               
                                                                                                                                         
        local_tmr_voter(325)  <=    (tmr_registers(0)(325) and tmr_registers(1)(325)) or                                                             
                            (tmr_registers(1)(325) and tmr_registers(2)(325)) or                                                             
                            (tmr_registers(0)(325) and tmr_registers(2)(325));                                                               
                                                                                                                                         
        local_tmr_voter(326)  <=    (tmr_registers(0)(326) and tmr_registers(1)(326)) or                                                             
                            (tmr_registers(1)(326) and tmr_registers(2)(326)) or                                                             
                            (tmr_registers(0)(326) and tmr_registers(2)(326));                                                               
                                                                                                                                         
        local_tmr_voter(327)  <=    (tmr_registers(0)(327) and tmr_registers(1)(327)) or                                                             
                            (tmr_registers(1)(327) and tmr_registers(2)(327)) or                                                             
                            (tmr_registers(0)(327) and tmr_registers(2)(327));                                                               
                                                                                                                                         
        local_tmr_voter(328)  <=    (tmr_registers(0)(328) and tmr_registers(1)(328)) or                                                             
                            (tmr_registers(1)(328) and tmr_registers(2)(328)) or                                                             
                            (tmr_registers(0)(328) and tmr_registers(2)(328));                                                               
                                                                                                                                         
        local_tmr_voter(329)  <=    (tmr_registers(0)(329) and tmr_registers(1)(329)) or                                                             
                            (tmr_registers(1)(329) and tmr_registers(2)(329)) or                                                             
                            (tmr_registers(0)(329) and tmr_registers(2)(329));                                                               
                                                                                                                                         
        local_tmr_voter(330)  <=    (tmr_registers(0)(330) and tmr_registers(1)(330)) or                                                             
                            (tmr_registers(1)(330) and tmr_registers(2)(330)) or                                                             
                            (tmr_registers(0)(330) and tmr_registers(2)(330));                                                               
                                                                                                                                         
        local_tmr_voter(331)  <=    (tmr_registers(0)(331) and tmr_registers(1)(331)) or                                                             
                            (tmr_registers(1)(331) and tmr_registers(2)(331)) or                                                             
                            (tmr_registers(0)(331) and tmr_registers(2)(331));                                                               
                                                                                                                                         
        local_tmr_voter(332)  <=    (tmr_registers(0)(332) and tmr_registers(1)(332)) or                                                             
                            (tmr_registers(1)(332) and tmr_registers(2)(332)) or                                                             
                            (tmr_registers(0)(332) and tmr_registers(2)(332));                                                               
                                                                                                                                         
        local_tmr_voter(333)  <=    (tmr_registers(0)(333) and tmr_registers(1)(333)) or                                                             
                            (tmr_registers(1)(333) and tmr_registers(2)(333)) or                                                             
                            (tmr_registers(0)(333) and tmr_registers(2)(333));                                                               
                                                                                                                                         
        local_tmr_voter(334)  <=    (tmr_registers(0)(334) and tmr_registers(1)(334)) or                                                             
                            (tmr_registers(1)(334) and tmr_registers(2)(334)) or                                                             
                            (tmr_registers(0)(334) and tmr_registers(2)(334));                                                               
                                                                                                                                         
        local_tmr_voter(335)  <=    (tmr_registers(0)(335) and tmr_registers(1)(335)) or                                                             
                            (tmr_registers(1)(335) and tmr_registers(2)(335)) or                                                             
                            (tmr_registers(0)(335) and tmr_registers(2)(335));                                                               
                                                                                                                                         
        local_tmr_voter(336)  <=    (tmr_registers(0)(336) and tmr_registers(1)(336)) or                                                             
                            (tmr_registers(1)(336) and tmr_registers(2)(336)) or                                                             
                            (tmr_registers(0)(336) and tmr_registers(2)(336));                                                               
                                                                                                                                         
        local_tmr_voter(337)  <=    (tmr_registers(0)(337) and tmr_registers(1)(337)) or                                                             
                            (tmr_registers(1)(337) and tmr_registers(2)(337)) or                                                             
                            (tmr_registers(0)(337) and tmr_registers(2)(337));                                                               
                                                                                                                                         
        local_tmr_voter(338)  <=    (tmr_registers(0)(338) and tmr_registers(1)(338)) or                                                             
                            (tmr_registers(1)(338) and tmr_registers(2)(338)) or                                                             
                            (tmr_registers(0)(338) and tmr_registers(2)(338));                                                               
                                                                                                                                         
        local_tmr_voter(339)  <=    (tmr_registers(0)(339) and tmr_registers(1)(339)) or                                                             
                            (tmr_registers(1)(339) and tmr_registers(2)(339)) or                                                             
                            (tmr_registers(0)(339) and tmr_registers(2)(339));                                                               
                                                                                                                                         
        local_tmr_voter(340)  <=    (tmr_registers(0)(340) and tmr_registers(1)(340)) or                                                             
                            (tmr_registers(1)(340) and tmr_registers(2)(340)) or                                                             
                            (tmr_registers(0)(340) and tmr_registers(2)(340));                                                               
                                                                                                                                         
        local_tmr_voter(341)  <=    (tmr_registers(0)(341) and tmr_registers(1)(341)) or                                                             
                            (tmr_registers(1)(341) and tmr_registers(2)(341)) or                                                             
                            (tmr_registers(0)(341) and tmr_registers(2)(341));                                                               
                                                                                                                                         
        local_tmr_voter(342)  <=    (tmr_registers(0)(342) and tmr_registers(1)(342)) or                                                             
                            (tmr_registers(1)(342) and tmr_registers(2)(342)) or                                                             
                            (tmr_registers(0)(342) and tmr_registers(2)(342));                                                               
                                                                                                                                         
        local_tmr_voter(343)  <=    (tmr_registers(0)(343) and tmr_registers(1)(343)) or                                                             
                            (tmr_registers(1)(343) and tmr_registers(2)(343)) or                                                             
                            (tmr_registers(0)(343) and tmr_registers(2)(343));                                                               
                                                                                                                                         
        local_tmr_voter(344)  <=    (tmr_registers(0)(344) and tmr_registers(1)(344)) or                                                             
                            (tmr_registers(1)(344) and tmr_registers(2)(344)) or                                                             
                            (tmr_registers(0)(344) and tmr_registers(2)(344));                                                               
                                                                                                                                         
        local_tmr_voter(345)  <=    (tmr_registers(0)(345) and tmr_registers(1)(345)) or                                                             
                            (tmr_registers(1)(345) and tmr_registers(2)(345)) or                                                             
                            (tmr_registers(0)(345) and tmr_registers(2)(345));                                                               
                                                                                                                                         
        local_tmr_voter(346)  <=    (tmr_registers(0)(346) and tmr_registers(1)(346)) or                                                             
                            (tmr_registers(1)(346) and tmr_registers(2)(346)) or                                                             
                            (tmr_registers(0)(346) and tmr_registers(2)(346));                                                               
                                                                                                                                         
        local_tmr_voter(347)  <=    (tmr_registers(0)(347) and tmr_registers(1)(347)) or                                                             
                            (tmr_registers(1)(347) and tmr_registers(2)(347)) or                                                             
                            (tmr_registers(0)(347) and tmr_registers(2)(347));                                                               
                                                                                                                                         
        local_tmr_voter(348)  <=    (tmr_registers(0)(348) and tmr_registers(1)(348)) or                                                             
                            (tmr_registers(1)(348) and tmr_registers(2)(348)) or                                                             
                            (tmr_registers(0)(348) and tmr_registers(2)(348));                                                               
                                                                                                                                         
        local_tmr_voter(349)  <=    (tmr_registers(0)(349) and tmr_registers(1)(349)) or                                                             
                            (tmr_registers(1)(349) and tmr_registers(2)(349)) or                                                             
                            (tmr_registers(0)(349) and tmr_registers(2)(349));                                                               
                                                                                                                                         
        local_tmr_voter(350)  <=    (tmr_registers(0)(350) and tmr_registers(1)(350)) or                                                             
                            (tmr_registers(1)(350) and tmr_registers(2)(350)) or                                                             
                            (tmr_registers(0)(350) and tmr_registers(2)(350));                                                               
                                                                                                                                         
        local_tmr_voter(351)  <=    (tmr_registers(0)(351) and tmr_registers(1)(351)) or                                                             
                            (tmr_registers(1)(351) and tmr_registers(2)(351)) or                                                             
                            (tmr_registers(0)(351) and tmr_registers(2)(351));                                                               
                                                                                                                                         
        local_tmr_voter(352)  <=    (tmr_registers(0)(352) and tmr_registers(1)(352)) or                                                             
                            (tmr_registers(1)(352) and tmr_registers(2)(352)) or                                                             
                            (tmr_registers(0)(352) and tmr_registers(2)(352));                                                               
                                                                                                                                         
        local_tmr_voter(353)  <=    (tmr_registers(0)(353) and tmr_registers(1)(353)) or                                                             
                            (tmr_registers(1)(353) and tmr_registers(2)(353)) or                                                             
                            (tmr_registers(0)(353) and tmr_registers(2)(353));                                                               
                                                                                                                                         
        local_tmr_voter(354)  <=    (tmr_registers(0)(354) and tmr_registers(1)(354)) or                                                             
                            (tmr_registers(1)(354) and tmr_registers(2)(354)) or                                                             
                            (tmr_registers(0)(354) and tmr_registers(2)(354));                                                               
                                                                                                                                         
        local_tmr_voter(355)  <=    (tmr_registers(0)(355) and tmr_registers(1)(355)) or                                                             
                            (tmr_registers(1)(355) and tmr_registers(2)(355)) or                                                             
                            (tmr_registers(0)(355) and tmr_registers(2)(355));                                                               
                                                                                                                                         
        local_tmr_voter(356)  <=    (tmr_registers(0)(356) and tmr_registers(1)(356)) or                                                             
                            (tmr_registers(1)(356) and tmr_registers(2)(356)) or                                                             
                            (tmr_registers(0)(356) and tmr_registers(2)(356));                                                               
                                                                                                                                         
        local_tmr_voter(357)  <=    (tmr_registers(0)(357) and tmr_registers(1)(357)) or                                                             
                            (tmr_registers(1)(357) and tmr_registers(2)(357)) or                                                             
                            (tmr_registers(0)(357) and tmr_registers(2)(357));                                                               
                                                                                                                                         
        local_tmr_voter(358)  <=    (tmr_registers(0)(358) and tmr_registers(1)(358)) or                                                             
                            (tmr_registers(1)(358) and tmr_registers(2)(358)) or                                                             
                            (tmr_registers(0)(358) and tmr_registers(2)(358));                                                               
                                                                                                                                         
        local_tmr_voter(359)  <=    (tmr_registers(0)(359) and tmr_registers(1)(359)) or                                                             
                            (tmr_registers(1)(359) and tmr_registers(2)(359)) or                                                             
                            (tmr_registers(0)(359) and tmr_registers(2)(359));                                                               
                                                                                                                                         
        local_tmr_voter(360)  <=    (tmr_registers(0)(360) and tmr_registers(1)(360)) or                                                             
                            (tmr_registers(1)(360) and tmr_registers(2)(360)) or                                                             
                            (tmr_registers(0)(360) and tmr_registers(2)(360));                                                               
                                                                                                                                         
        local_tmr_voter(361)  <=    (tmr_registers(0)(361) and tmr_registers(1)(361)) or                                                             
                            (tmr_registers(1)(361) and tmr_registers(2)(361)) or                                                             
                            (tmr_registers(0)(361) and tmr_registers(2)(361));                                                               
                                                                                                                                         
        local_tmr_voter(362)  <=    (tmr_registers(0)(362) and tmr_registers(1)(362)) or                                                             
                            (tmr_registers(1)(362) and tmr_registers(2)(362)) or                                                             
                            (tmr_registers(0)(362) and tmr_registers(2)(362));                                                               
                                                                                                                                         
        local_tmr_voter(363)  <=    (tmr_registers(0)(363) and tmr_registers(1)(363)) or                                                             
                            (tmr_registers(1)(363) and tmr_registers(2)(363)) or                                                             
                            (tmr_registers(0)(363) and tmr_registers(2)(363));                                                               
                                                                                                                                         
        local_tmr_voter(364)  <=    (tmr_registers(0)(364) and tmr_registers(1)(364)) or                                                             
                            (tmr_registers(1)(364) and tmr_registers(2)(364)) or                                                             
                            (tmr_registers(0)(364) and tmr_registers(2)(364));                                                               
                                                                                                                                         
        local_tmr_voter(365)  <=    (tmr_registers(0)(365) and tmr_registers(1)(365)) or                                                             
                            (tmr_registers(1)(365) and tmr_registers(2)(365)) or                                                             
                            (tmr_registers(0)(365) and tmr_registers(2)(365));                                                               
                                                                                                                                         
        local_tmr_voter(366)  <=    (tmr_registers(0)(366) and tmr_registers(1)(366)) or                                                             
                            (tmr_registers(1)(366) and tmr_registers(2)(366)) or                                                             
                            (tmr_registers(0)(366) and tmr_registers(2)(366));                                                               
                                                                                                                                         
        local_tmr_voter(367)  <=    (tmr_registers(0)(367) and tmr_registers(1)(367)) or                                                             
                            (tmr_registers(1)(367) and tmr_registers(2)(367)) or                                                             
                            (tmr_registers(0)(367) and tmr_registers(2)(367));                                                               
                                                                                                                                         
        local_tmr_voter(368)  <=    (tmr_registers(0)(368) and tmr_registers(1)(368)) or                                                             
                            (tmr_registers(1)(368) and tmr_registers(2)(368)) or                                                             
                            (tmr_registers(0)(368) and tmr_registers(2)(368));                                                               
                                                                                                                                         
        local_tmr_voter(369)  <=    (tmr_registers(0)(369) and tmr_registers(1)(369)) or                                                             
                            (tmr_registers(1)(369) and tmr_registers(2)(369)) or                                                             
                            (tmr_registers(0)(369) and tmr_registers(2)(369));                                                               
                                                                                                                                         
        local_tmr_voter(370)  <=    (tmr_registers(0)(370) and tmr_registers(1)(370)) or                                                             
                            (tmr_registers(1)(370) and tmr_registers(2)(370)) or                                                             
                            (tmr_registers(0)(370) and tmr_registers(2)(370));                                                               
                                                                                                                                         
        local_tmr_voter(371)  <=    (tmr_registers(0)(371) and tmr_registers(1)(371)) or                                                             
                            (tmr_registers(1)(371) and tmr_registers(2)(371)) or                                                             
                            (tmr_registers(0)(371) and tmr_registers(2)(371));                                                               
                                                                                                                                         
        local_tmr_voter(372)  <=    (tmr_registers(0)(372) and tmr_registers(1)(372)) or                                                             
                            (tmr_registers(1)(372) and tmr_registers(2)(372)) or                                                             
                            (tmr_registers(0)(372) and tmr_registers(2)(372));                                                               
                                                                                                                                         
        local_tmr_voter(373)  <=    (tmr_registers(0)(373) and tmr_registers(1)(373)) or                                                             
                            (tmr_registers(1)(373) and tmr_registers(2)(373)) or                                                             
                            (tmr_registers(0)(373) and tmr_registers(2)(373));                                                               
                                                                                                                                         
        local_tmr_voter(374)  <=    (tmr_registers(0)(374) and tmr_registers(1)(374)) or                                                             
                            (tmr_registers(1)(374) and tmr_registers(2)(374)) or                                                             
                            (tmr_registers(0)(374) and tmr_registers(2)(374));                                                               
                                                                                                                                         
        local_tmr_voter(375)  <=    (tmr_registers(0)(375) and tmr_registers(1)(375)) or                                                             
                            (tmr_registers(1)(375) and tmr_registers(2)(375)) or                                                             
                            (tmr_registers(0)(375) and tmr_registers(2)(375));                                                               
                                                                                                                                         
        local_tmr_voter(376)  <=    (tmr_registers(0)(376) and tmr_registers(1)(376)) or                                                             
                            (tmr_registers(1)(376) and tmr_registers(2)(376)) or                                                             
                            (tmr_registers(0)(376) and tmr_registers(2)(376));                                                               
                                                                                                                                         
        local_tmr_voter(377)  <=    (tmr_registers(0)(377) and tmr_registers(1)(377)) or                                                             
                            (tmr_registers(1)(377) and tmr_registers(2)(377)) or                                                             
                            (tmr_registers(0)(377) and tmr_registers(2)(377));                                                               
                                                                                                                                         
        local_tmr_voter(378)  <=    (tmr_registers(0)(378) and tmr_registers(1)(378)) or                                                             
                            (tmr_registers(1)(378) and tmr_registers(2)(378)) or                                                             
                            (tmr_registers(0)(378) and tmr_registers(2)(378));                                                               
                                                                                                                                         
        local_tmr_voter(379)  <=    (tmr_registers(0)(379) and tmr_registers(1)(379)) or                                                             
                            (tmr_registers(1)(379) and tmr_registers(2)(379)) or                                                             
                            (tmr_registers(0)(379) and tmr_registers(2)(379));                                                               
                                                                                                                                         
        local_tmr_voter(380)  <=    (tmr_registers(0)(380) and tmr_registers(1)(380)) or                                                             
                            (tmr_registers(1)(380) and tmr_registers(2)(380)) or                                                             
                            (tmr_registers(0)(380) and tmr_registers(2)(380));                                                               
                                                                                                                                         
        local_tmr_voter(381)  <=    (tmr_registers(0)(381) and tmr_registers(1)(381)) or                                                             
                            (tmr_registers(1)(381) and tmr_registers(2)(381)) or                                                             
                            (tmr_registers(0)(381) and tmr_registers(2)(381));                                                               
                                                                                                                                         
        local_tmr_voter(382)  <=    (tmr_registers(0)(382) and tmr_registers(1)(382)) or                                                             
                            (tmr_registers(1)(382) and tmr_registers(2)(382)) or                                                             
                            (tmr_registers(0)(382) and tmr_registers(2)(382));                                                               
                                                                                                                                         
        local_tmr_voter(383)  <=    (tmr_registers(0)(383) and tmr_registers(1)(383)) or                                                             
                            (tmr_registers(1)(383) and tmr_registers(2)(383)) or                                                             
                            (tmr_registers(0)(383) and tmr_registers(2)(383));                                                               
                                                                                                                                         
        local_tmr_voter(384)  <=    (tmr_registers(0)(384) and tmr_registers(1)(384)) or                                                             
                            (tmr_registers(1)(384) and tmr_registers(2)(384)) or                                                             
                            (tmr_registers(0)(384) and tmr_registers(2)(384));                                                               
                                                                                                                                         
        local_tmr_voter(385)  <=    (tmr_registers(0)(385) and tmr_registers(1)(385)) or                                                             
                            (tmr_registers(1)(385) and tmr_registers(2)(385)) or                                                             
                            (tmr_registers(0)(385) and tmr_registers(2)(385));                                                               
                                                                                                                                         
        local_tmr_voter(386)  <=    (tmr_registers(0)(386) and tmr_registers(1)(386)) or                                                             
                            (tmr_registers(1)(386) and tmr_registers(2)(386)) or                                                             
                            (tmr_registers(0)(386) and tmr_registers(2)(386));                                                               
                                                                                                                                         
        local_tmr_voter(387)  <=    (tmr_registers(0)(387) and tmr_registers(1)(387)) or                                                             
                            (tmr_registers(1)(387) and tmr_registers(2)(387)) or                                                             
                            (tmr_registers(0)(387) and tmr_registers(2)(387));                                                               
                                                                                                                                         
        local_tmr_voter(388)  <=    (tmr_registers(0)(388) and tmr_registers(1)(388)) or                                                             
                            (tmr_registers(1)(388) and tmr_registers(2)(388)) or                                                             
                            (tmr_registers(0)(388) and tmr_registers(2)(388));                                                               
                                                                                                                                         
        local_tmr_voter(389)  <=    (tmr_registers(0)(389) and tmr_registers(1)(389)) or                                                             
                            (tmr_registers(1)(389) and tmr_registers(2)(389)) or                                                             
                            (tmr_registers(0)(389) and tmr_registers(2)(389));                                                               
                                                                                                                                         
        local_tmr_voter(390)  <=    (tmr_registers(0)(390) and tmr_registers(1)(390)) or                                                             
                            (tmr_registers(1)(390) and tmr_registers(2)(390)) or                                                             
                            (tmr_registers(0)(390) and tmr_registers(2)(390));                                                               
                                                                                                                                         
        local_tmr_voter(391)  <=    (tmr_registers(0)(391) and tmr_registers(1)(391)) or                                                             
                            (tmr_registers(1)(391) and tmr_registers(2)(391)) or                                                             
                            (tmr_registers(0)(391) and tmr_registers(2)(391));                                                               
                                                                                                                                         
        local_tmr_voter(392)  <=    (tmr_registers(0)(392) and tmr_registers(1)(392)) or                                                             
                            (tmr_registers(1)(392) and tmr_registers(2)(392)) or                                                             
                            (tmr_registers(0)(392) and tmr_registers(2)(392));                                                               
                                                                                                                                         
        local_tmr_voter(393)  <=    (tmr_registers(0)(393) and tmr_registers(1)(393)) or                                                             
                            (tmr_registers(1)(393) and tmr_registers(2)(393)) or                                                             
                            (tmr_registers(0)(393) and tmr_registers(2)(393));                                                               
                                                                                                                                         
        local_tmr_voter(394)  <=    (tmr_registers(0)(394) and tmr_registers(1)(394)) or                                                             
                            (tmr_registers(1)(394) and tmr_registers(2)(394)) or                                                             
                            (tmr_registers(0)(394) and tmr_registers(2)(394));                                                               
                                                                                                                                         
        local_tmr_voter(395)  <=    (tmr_registers(0)(395) and tmr_registers(1)(395)) or                                                             
                            (tmr_registers(1)(395) and tmr_registers(2)(395)) or                                                             
                            (tmr_registers(0)(395) and tmr_registers(2)(395));                                                               
                                                                                                                                         
        local_tmr_voter(396)  <=    (tmr_registers(0)(396) and tmr_registers(1)(396)) or                                                             
                            (tmr_registers(1)(396) and tmr_registers(2)(396)) or                                                             
                            (tmr_registers(0)(396) and tmr_registers(2)(396));                                                               
                                                                                                                                         
        local_tmr_voter(397)  <=    (tmr_registers(0)(397) and tmr_registers(1)(397)) or                                                             
                            (tmr_registers(1)(397) and tmr_registers(2)(397)) or                                                             
                            (tmr_registers(0)(397) and tmr_registers(2)(397));                                                               
                                                                                                                                         
        local_tmr_voter(398)  <=    (tmr_registers(0)(398) and tmr_registers(1)(398)) or                                                             
                            (tmr_registers(1)(398) and tmr_registers(2)(398)) or                                                             
                            (tmr_registers(0)(398) and tmr_registers(2)(398));                                                               
                                                                                                                                         
        local_tmr_voter(399)  <=    (tmr_registers(0)(399) and tmr_registers(1)(399)) or                                                             
                            (tmr_registers(1)(399) and tmr_registers(2)(399)) or                                                             
                            (tmr_registers(0)(399) and tmr_registers(2)(399));                                                               
                                                                                                                                         
        local_tmr_voter(400)  <=    (tmr_registers(0)(400) and tmr_registers(1)(400)) or                                                             
                            (tmr_registers(1)(400) and tmr_registers(2)(400)) or                                                             
                            (tmr_registers(0)(400) and tmr_registers(2)(400));                                                               
                                                                                                                                         
        local_tmr_voter(401)  <=    (tmr_registers(0)(401) and tmr_registers(1)(401)) or                                                             
                            (tmr_registers(1)(401) and tmr_registers(2)(401)) or                                                             
                            (tmr_registers(0)(401) and tmr_registers(2)(401));                                                               
                                                                                                                                         
        local_tmr_voter(402)  <=    (tmr_registers(0)(402) and tmr_registers(1)(402)) or                                                             
                            (tmr_registers(1)(402) and tmr_registers(2)(402)) or                                                             
                            (tmr_registers(0)(402) and tmr_registers(2)(402));                                                               
                                                                                                                                         
        local_tmr_voter(403)  <=    (tmr_registers(0)(403) and tmr_registers(1)(403)) or                                                             
                            (tmr_registers(1)(403) and tmr_registers(2)(403)) or                                                             
                            (tmr_registers(0)(403) and tmr_registers(2)(403));                                                               
                                                                                                                                         
        local_tmr_voter(404)  <=    (tmr_registers(0)(404) and tmr_registers(1)(404)) or                                                             
                            (tmr_registers(1)(404) and tmr_registers(2)(404)) or                                                             
                            (tmr_registers(0)(404) and tmr_registers(2)(404));                                                               
                                                                                                                                         
        local_tmr_voter(405)  <=    (tmr_registers(0)(405) and tmr_registers(1)(405)) or                                                             
                            (tmr_registers(1)(405) and tmr_registers(2)(405)) or                                                             
                            (tmr_registers(0)(405) and tmr_registers(2)(405));                                                               
                                                                                                                                         
        local_tmr_voter(406)  <=    (tmr_registers(0)(406) and tmr_registers(1)(406)) or                                                             
                            (tmr_registers(1)(406) and tmr_registers(2)(406)) or                                                             
                            (tmr_registers(0)(406) and tmr_registers(2)(406));                                                               
                                                                                                                                         
        local_tmr_voter(407)  <=    (tmr_registers(0)(407) and tmr_registers(1)(407)) or                                                             
                            (tmr_registers(1)(407) and tmr_registers(2)(407)) or                                                             
                            (tmr_registers(0)(407) and tmr_registers(2)(407));                                                               
                                                                                                                                         
        local_tmr_voter(408)  <=    (tmr_registers(0)(408) and tmr_registers(1)(408)) or                                                             
                            (tmr_registers(1)(408) and tmr_registers(2)(408)) or                                                             
                            (tmr_registers(0)(408) and tmr_registers(2)(408));                                                               
                                                                                                                                         
        local_tmr_voter(409)  <=    (tmr_registers(0)(409) and tmr_registers(1)(409)) or                                                             
                            (tmr_registers(1)(409) and tmr_registers(2)(409)) or                                                             
                            (tmr_registers(0)(409) and tmr_registers(2)(409));                                                               
                                                                                                                                         
        local_tmr_voter(410)  <=    (tmr_registers(0)(410) and tmr_registers(1)(410)) or                                                             
                            (tmr_registers(1)(410) and tmr_registers(2)(410)) or                                                             
                            (tmr_registers(0)(410) and tmr_registers(2)(410));                                                               
                                                                                                                                         
        local_tmr_voter(411)  <=    (tmr_registers(0)(411) and tmr_registers(1)(411)) or                                                             
                            (tmr_registers(1)(411) and tmr_registers(2)(411)) or                                                             
                            (tmr_registers(0)(411) and tmr_registers(2)(411));                                                               
                                                                                                                                         
        local_tmr_voter(412)  <=    (tmr_registers(0)(412) and tmr_registers(1)(412)) or                                                             
                            (tmr_registers(1)(412) and tmr_registers(2)(412)) or                                                             
                            (tmr_registers(0)(412) and tmr_registers(2)(412));                                                               
                                                                                                                                         
        local_tmr_voter(413)  <=    (tmr_registers(0)(413) and tmr_registers(1)(413)) or                                                             
                            (tmr_registers(1)(413) and tmr_registers(2)(413)) or                                                             
                            (tmr_registers(0)(413) and tmr_registers(2)(413));                                                               
                                                                                                                                         
        local_tmr_voter(414)  <=    (tmr_registers(0)(414) and tmr_registers(1)(414)) or                                                             
                            (tmr_registers(1)(414) and tmr_registers(2)(414)) or                                                             
                            (tmr_registers(0)(414) and tmr_registers(2)(414));                                                               
                                                                                                                                         
        local_tmr_voter(415)  <=    (tmr_registers(0)(415) and tmr_registers(1)(415)) or                                                             
                            (tmr_registers(1)(415) and tmr_registers(2)(415)) or                                                             
                            (tmr_registers(0)(415) and tmr_registers(2)(415));                                                               
                                                                                                                                         
        local_tmr_voter(416)  <=    (tmr_registers(0)(416) and tmr_registers(1)(416)) or                                                             
                            (tmr_registers(1)(416) and tmr_registers(2)(416)) or                                                             
                            (tmr_registers(0)(416) and tmr_registers(2)(416));                                                               
                                                                                                                                         
        local_tmr_voter(417)  <=    (tmr_registers(0)(417) and tmr_registers(1)(417)) or                                                             
                            (tmr_registers(1)(417) and tmr_registers(2)(417)) or                                                             
                            (tmr_registers(0)(417) and tmr_registers(2)(417));                                                               
                                                                                                                                         
        local_tmr_voter(418)  <=    (tmr_registers(0)(418) and tmr_registers(1)(418)) or                                                             
                            (tmr_registers(1)(418) and tmr_registers(2)(418)) or                                                             
                            (tmr_registers(0)(418) and tmr_registers(2)(418));                                                               
                                                                                                                                         
        local_tmr_voter(419)  <=    (tmr_registers(0)(419) and tmr_registers(1)(419)) or                                                             
                            (tmr_registers(1)(419) and tmr_registers(2)(419)) or                                                             
                            (tmr_registers(0)(419) and tmr_registers(2)(419));                                                               
                                                                                                                                         
        local_tmr_voter(420)  <=    (tmr_registers(0)(420) and tmr_registers(1)(420)) or                                                             
                            (tmr_registers(1)(420) and tmr_registers(2)(420)) or                                                             
                            (tmr_registers(0)(420) and tmr_registers(2)(420));                                                               
                                                                                                                                         
        local_tmr_voter(421)  <=    (tmr_registers(0)(421) and tmr_registers(1)(421)) or                                                             
                            (tmr_registers(1)(421) and tmr_registers(2)(421)) or                                                             
                            (tmr_registers(0)(421) and tmr_registers(2)(421));                                                               
                                                                                                                                         
        local_tmr_voter(422)  <=    (tmr_registers(0)(422) and tmr_registers(1)(422)) or                                                             
                            (tmr_registers(1)(422) and tmr_registers(2)(422)) or                                                             
                            (tmr_registers(0)(422) and tmr_registers(2)(422));                                                               
                                                                                                                                         
        local_tmr_voter(423)  <=    (tmr_registers(0)(423) and tmr_registers(1)(423)) or                                                             
                            (tmr_registers(1)(423) and tmr_registers(2)(423)) or                                                             
                            (tmr_registers(0)(423) and tmr_registers(2)(423));                                                               
                                                                                                                                         
        local_tmr_voter(424)  <=    (tmr_registers(0)(424) and tmr_registers(1)(424)) or                                                             
                            (tmr_registers(1)(424) and tmr_registers(2)(424)) or                                                             
                            (tmr_registers(0)(424) and tmr_registers(2)(424));                                                               
                                                                                                                                         
        local_tmr_voter(425)  <=    (tmr_registers(0)(425) and tmr_registers(1)(425)) or                                                             
                            (tmr_registers(1)(425) and tmr_registers(2)(425)) or                                                             
                            (tmr_registers(0)(425) and tmr_registers(2)(425));                                                               
                                                                                                                                         
        local_tmr_voter(426)  <=    (tmr_registers(0)(426) and tmr_registers(1)(426)) or                                                             
                            (tmr_registers(1)(426) and tmr_registers(2)(426)) or                                                             
                            (tmr_registers(0)(426) and tmr_registers(2)(426));                                                               
                                                                                                                                         
        local_tmr_voter(427)  <=    (tmr_registers(0)(427) and tmr_registers(1)(427)) or                                                             
                            (tmr_registers(1)(427) and tmr_registers(2)(427)) or                                                             
                            (tmr_registers(0)(427) and tmr_registers(2)(427));                                                               
                                                                                                                                         
        local_tmr_voter(428)  <=    (tmr_registers(0)(428) and tmr_registers(1)(428)) or                                                             
                            (tmr_registers(1)(428) and tmr_registers(2)(428)) or                                                             
                            (tmr_registers(0)(428) and tmr_registers(2)(428));                                                               
                                                                                                                                         
        local_tmr_voter(429)  <=    (tmr_registers(0)(429) and tmr_registers(1)(429)) or                                                             
                            (tmr_registers(1)(429) and tmr_registers(2)(429)) or                                                             
                            (tmr_registers(0)(429) and tmr_registers(2)(429));                                                               
                                                                                                                                         
        local_tmr_voter(430)  <=    (tmr_registers(0)(430) and tmr_registers(1)(430)) or                                                             
                            (tmr_registers(1)(430) and tmr_registers(2)(430)) or                                                             
                            (tmr_registers(0)(430) and tmr_registers(2)(430));                                                               
                                                                                                                                         
        local_tmr_voter(431)  <=    (tmr_registers(0)(431) and tmr_registers(1)(431)) or                                                             
                            (tmr_registers(1)(431) and tmr_registers(2)(431)) or                                                             
                            (tmr_registers(0)(431) and tmr_registers(2)(431));                                                               
                                                                                                                                         
        local_tmr_voter(432)  <=    (tmr_registers(0)(432) and tmr_registers(1)(432)) or                                                             
                            (tmr_registers(1)(432) and tmr_registers(2)(432)) or                                                             
                            (tmr_registers(0)(432) and tmr_registers(2)(432));                                                               
                                                                                                                                         
        local_tmr_voter(433)  <=    (tmr_registers(0)(433) and tmr_registers(1)(433)) or                                                             
                            (tmr_registers(1)(433) and tmr_registers(2)(433)) or                                                             
                            (tmr_registers(0)(433) and tmr_registers(2)(433));                                                               
                                                                                                                                         
        local_tmr_voter(434)  <=    (tmr_registers(0)(434) and tmr_registers(1)(434)) or                                                             
                            (tmr_registers(1)(434) and tmr_registers(2)(434)) or                                                             
                            (tmr_registers(0)(434) and tmr_registers(2)(434));                                                               
                                                                                                                                         
        local_tmr_voter(435)  <=    (tmr_registers(0)(435) and tmr_registers(1)(435)) or                                                             
                            (tmr_registers(1)(435) and tmr_registers(2)(435)) or                                                             
                            (tmr_registers(0)(435) and tmr_registers(2)(435));                                                               
                                                                                                                                         
        local_tmr_voter(436)  <=    (tmr_registers(0)(436) and tmr_registers(1)(436)) or                                                             
                            (tmr_registers(1)(436) and tmr_registers(2)(436)) or                                                             
                            (tmr_registers(0)(436) and tmr_registers(2)(436));                                                               
                                                                                                                                         
        local_tmr_voter(437)  <=    (tmr_registers(0)(437) and tmr_registers(1)(437)) or                                                             
                            (tmr_registers(1)(437) and tmr_registers(2)(437)) or                                                             
                            (tmr_registers(0)(437) and tmr_registers(2)(437));                                                               
                                                                                                                                         
        local_tmr_voter(438)  <=    (tmr_registers(0)(438) and tmr_registers(1)(438)) or                                                             
                            (tmr_registers(1)(438) and tmr_registers(2)(438)) or                                                             
                            (tmr_registers(0)(438) and tmr_registers(2)(438));                                                               
                                                                                                                                         
        local_tmr_voter(439)  <=    (tmr_registers(0)(439) and tmr_registers(1)(439)) or                                                             
                            (tmr_registers(1)(439) and tmr_registers(2)(439)) or                                                             
                            (tmr_registers(0)(439) and tmr_registers(2)(439));                                                               
                                                                                                                                         
        local_tmr_voter(440)  <=    (tmr_registers(0)(440) and tmr_registers(1)(440)) or                                                             
                            (tmr_registers(1)(440) and tmr_registers(2)(440)) or                                                             
                            (tmr_registers(0)(440) and tmr_registers(2)(440));                                                               
                                                                                                                                         
        local_tmr_voter(441)  <=    (tmr_registers(0)(441) and tmr_registers(1)(441)) or                                                             
                            (tmr_registers(1)(441) and tmr_registers(2)(441)) or                                                             
                            (tmr_registers(0)(441) and tmr_registers(2)(441));                                                               
                                                                                                                                         
        local_tmr_voter(442)  <=    (tmr_registers(0)(442) and tmr_registers(1)(442)) or                                                             
                            (tmr_registers(1)(442) and tmr_registers(2)(442)) or                                                             
                            (tmr_registers(0)(442) and tmr_registers(2)(442));                                                               
                                                                                                                                         
        local_tmr_voter(443)  <=    (tmr_registers(0)(443) and tmr_registers(1)(443)) or                                                             
                            (tmr_registers(1)(443) and tmr_registers(2)(443)) or                                                             
                            (tmr_registers(0)(443) and tmr_registers(2)(443));                                                               
                                                                                                                                         
        local_tmr_voter(444)  <=    (tmr_registers(0)(444) and tmr_registers(1)(444)) or                                                             
                            (tmr_registers(1)(444) and tmr_registers(2)(444)) or                                                             
                            (tmr_registers(0)(444) and tmr_registers(2)(444));                                                               
                                                                                                                                         
        local_tmr_voter(445)  <=    (tmr_registers(0)(445) and tmr_registers(1)(445)) or                                                             
                            (tmr_registers(1)(445) and tmr_registers(2)(445)) or                                                             
                            (tmr_registers(0)(445) and tmr_registers(2)(445));                                                               
                                                                                                                                         
        local_tmr_voter(446)  <=    (tmr_registers(0)(446) and tmr_registers(1)(446)) or                                                             
                            (tmr_registers(1)(446) and tmr_registers(2)(446)) or                                                             
                            (tmr_registers(0)(446) and tmr_registers(2)(446));                                                               
                                                                                                                                         
        local_tmr_voter(447)  <=    (tmr_registers(0)(447) and tmr_registers(1)(447)) or                                                             
                            (tmr_registers(1)(447) and tmr_registers(2)(447)) or                                                             
                            (tmr_registers(0)(447) and tmr_registers(2)(447));                                                               
                                                                                                                                         
        local_tmr_voter(448)  <=    (tmr_registers(0)(448) and tmr_registers(1)(448)) or                                                             
                            (tmr_registers(1)(448) and tmr_registers(2)(448)) or                                                             
                            (tmr_registers(0)(448) and tmr_registers(2)(448));                                                               
                                                                                                                                         
        local_tmr_voter(449)  <=    (tmr_registers(0)(449) and tmr_registers(1)(449)) or                                                             
                            (tmr_registers(1)(449) and tmr_registers(2)(449)) or                                                             
                            (tmr_registers(0)(449) and tmr_registers(2)(449));                                                               
                                                                                                                                         
        local_tmr_voter(450)  <=    (tmr_registers(0)(450) and tmr_registers(1)(450)) or                                                             
                            (tmr_registers(1)(450) and tmr_registers(2)(450)) or                                                             
                            (tmr_registers(0)(450) and tmr_registers(2)(450));                                                               
                                                                                                                                         
        local_tmr_voter(451)  <=    (tmr_registers(0)(451) and tmr_registers(1)(451)) or                                                             
                            (tmr_registers(1)(451) and tmr_registers(2)(451)) or                                                             
                            (tmr_registers(0)(451) and tmr_registers(2)(451));                                                               
                                                                                                                                         
        local_tmr_voter(452)  <=    (tmr_registers(0)(452) and tmr_registers(1)(452)) or                                                             
                            (tmr_registers(1)(452) and tmr_registers(2)(452)) or                                                             
                            (tmr_registers(0)(452) and tmr_registers(2)(452));                                                               
                                                                                                                                         
        local_tmr_voter(453)  <=    (tmr_registers(0)(453) and tmr_registers(1)(453)) or                                                             
                            (tmr_registers(1)(453) and tmr_registers(2)(453)) or                                                             
                            (tmr_registers(0)(453) and tmr_registers(2)(453));                                                               
                                                                                                                                         
        local_tmr_voter(454)  <=    (tmr_registers(0)(454) and tmr_registers(1)(454)) or                                                             
                            (tmr_registers(1)(454) and tmr_registers(2)(454)) or                                                             
                            (tmr_registers(0)(454) and tmr_registers(2)(454));                                                               
                                                                                                                                         
        local_tmr_voter(455)  <=    (tmr_registers(0)(455) and tmr_registers(1)(455)) or                                                             
                            (tmr_registers(1)(455) and tmr_registers(2)(455)) or                                                             
                            (tmr_registers(0)(455) and tmr_registers(2)(455));                                                               
                                                                                                                                         
        local_tmr_voter(456)  <=    (tmr_registers(0)(456) and tmr_registers(1)(456)) or                                                             
                            (tmr_registers(1)(456) and tmr_registers(2)(456)) or                                                             
                            (tmr_registers(0)(456) and tmr_registers(2)(456));                                                               
                                                                                                                                         
        local_tmr_voter(457)  <=    (tmr_registers(0)(457) and tmr_registers(1)(457)) or                                                             
                            (tmr_registers(1)(457) and tmr_registers(2)(457)) or                                                             
                            (tmr_registers(0)(457) and tmr_registers(2)(457));                                                               
                                                                                                                                         
        local_tmr_voter(458)  <=    (tmr_registers(0)(458) and tmr_registers(1)(458)) or                                                             
                            (tmr_registers(1)(458) and tmr_registers(2)(458)) or                                                             
                            (tmr_registers(0)(458) and tmr_registers(2)(458));                                                               
                                                                                                                                         
        local_tmr_voter(459)  <=    (tmr_registers(0)(459) and tmr_registers(1)(459)) or                                                             
                            (tmr_registers(1)(459) and tmr_registers(2)(459)) or                                                             
                            (tmr_registers(0)(459) and tmr_registers(2)(459));                                                               
                                                                                                                                         
        local_tmr_voter(460)  <=    (tmr_registers(0)(460) and tmr_registers(1)(460)) or                                                             
                            (tmr_registers(1)(460) and tmr_registers(2)(460)) or                                                             
                            (tmr_registers(0)(460) and tmr_registers(2)(460));                                                               
                                                                                                                                         
        local_tmr_voter(461)  <=    (tmr_registers(0)(461) and tmr_registers(1)(461)) or                                                             
                            (tmr_registers(1)(461) and tmr_registers(2)(461)) or                                                             
                            (tmr_registers(0)(461) and tmr_registers(2)(461));                                                               
                                                                                                                                         
        local_tmr_voter(462)  <=    (tmr_registers(0)(462) and tmr_registers(1)(462)) or                                                             
                            (tmr_registers(1)(462) and tmr_registers(2)(462)) or                                                             
                            (tmr_registers(0)(462) and tmr_registers(2)(462));                                                               
                                                                                                                                         
        local_tmr_voter(463)  <=    (tmr_registers(0)(463) and tmr_registers(1)(463)) or                                                             
                            (tmr_registers(1)(463) and tmr_registers(2)(463)) or                                                             
                            (tmr_registers(0)(463) and tmr_registers(2)(463));                                                               
                                                                                                                                         
        local_tmr_voter(464)  <=    (tmr_registers(0)(464) and tmr_registers(1)(464)) or                                                             
                            (tmr_registers(1)(464) and tmr_registers(2)(464)) or                                                             
                            (tmr_registers(0)(464) and tmr_registers(2)(464));                                                               
                                                                                                                                         
        local_tmr_voter(465)  <=    (tmr_registers(0)(465) and tmr_registers(1)(465)) or                                                             
                            (tmr_registers(1)(465) and tmr_registers(2)(465)) or                                                             
                            (tmr_registers(0)(465) and tmr_registers(2)(465));                                                               
                                                                                                                                         
        local_tmr_voter(466)  <=    (tmr_registers(0)(466) and tmr_registers(1)(466)) or                                                             
                            (tmr_registers(1)(466) and tmr_registers(2)(466)) or                                                             
                            (tmr_registers(0)(466) and tmr_registers(2)(466));                                                               
                                                                                                                                         
        local_tmr_voter(467)  <=    (tmr_registers(0)(467) and tmr_registers(1)(467)) or                                                             
                            (tmr_registers(1)(467) and tmr_registers(2)(467)) or                                                             
                            (tmr_registers(0)(467) and tmr_registers(2)(467));                                                               
                                                                                                                                         
        local_tmr_voter(468)  <=    (tmr_registers(0)(468) and tmr_registers(1)(468)) or                                                             
                            (tmr_registers(1)(468) and tmr_registers(2)(468)) or                                                             
                            (tmr_registers(0)(468) and tmr_registers(2)(468));                                                               
                                                                                                                                         
        local_tmr_voter(469)  <=    (tmr_registers(0)(469) and tmr_registers(1)(469)) or                                                             
                            (tmr_registers(1)(469) and tmr_registers(2)(469)) or                                                             
                            (tmr_registers(0)(469) and tmr_registers(2)(469));                                                               
                                                                                                                                         
        local_tmr_voter(470)  <=    (tmr_registers(0)(470) and tmr_registers(1)(470)) or                                                             
                            (tmr_registers(1)(470) and tmr_registers(2)(470)) or                                                             
                            (tmr_registers(0)(470) and tmr_registers(2)(470));                                                               
                                                                                                                                         
        local_tmr_voter(471)  <=    (tmr_registers(0)(471) and tmr_registers(1)(471)) or                                                             
                            (tmr_registers(1)(471) and tmr_registers(2)(471)) or                                                             
                            (tmr_registers(0)(471) and tmr_registers(2)(471));                                                               
                                                                                                                                         
        local_tmr_voter(472)  <=    (tmr_registers(0)(472) and tmr_registers(1)(472)) or                                                             
                            (tmr_registers(1)(472) and tmr_registers(2)(472)) or                                                             
                            (tmr_registers(0)(472) and tmr_registers(2)(472));                                                               
                                                                                                                                         
        local_tmr_voter(473)  <=    (tmr_registers(0)(473) and tmr_registers(1)(473)) or                                                             
                            (tmr_registers(1)(473) and tmr_registers(2)(473)) or                                                             
                            (tmr_registers(0)(473) and tmr_registers(2)(473));                                                               
                                                                                                                                         
        local_tmr_voter(474)  <=    (tmr_registers(0)(474) and tmr_registers(1)(474)) or                                                             
                            (tmr_registers(1)(474) and tmr_registers(2)(474)) or                                                             
                            (tmr_registers(0)(474) and tmr_registers(2)(474));                                                               
                                                                                                                                         
        local_tmr_voter(475)  <=    (tmr_registers(0)(475) and tmr_registers(1)(475)) or                                                             
                            (tmr_registers(1)(475) and tmr_registers(2)(475)) or                                                             
                            (tmr_registers(0)(475) and tmr_registers(2)(475));                                                               
                                                                                                                                         
        local_tmr_voter(476)  <=    (tmr_registers(0)(476) and tmr_registers(1)(476)) or                                                             
                            (tmr_registers(1)(476) and tmr_registers(2)(476)) or                                                             
                            (tmr_registers(0)(476) and tmr_registers(2)(476));                                                               
                                                                                                                                         
        local_tmr_voter(477)  <=    (tmr_registers(0)(477) and tmr_registers(1)(477)) or                                                             
                            (tmr_registers(1)(477) and tmr_registers(2)(477)) or                                                             
                            (tmr_registers(0)(477) and tmr_registers(2)(477));                                                               
                                                                                                                                         
        local_tmr_voter(478)  <=    (tmr_registers(0)(478) and tmr_registers(1)(478)) or                                                             
                            (tmr_registers(1)(478) and tmr_registers(2)(478)) or                                                             
                            (tmr_registers(0)(478) and tmr_registers(2)(478));                                                               
                                                                                                                                         
        local_tmr_voter(479)  <=    (tmr_registers(0)(479) and tmr_registers(1)(479)) or                                                             
                            (tmr_registers(1)(479) and tmr_registers(2)(479)) or                                                             
                            (tmr_registers(0)(479) and tmr_registers(2)(479));                                                               
                                                                                                                                         
        local_tmr_voter(480)  <=    (tmr_registers(0)(480) and tmr_registers(1)(480)) or                                                             
                            (tmr_registers(1)(480) and tmr_registers(2)(480)) or                                                             
                            (tmr_registers(0)(480) and tmr_registers(2)(480));                                                               
                                                                                                                                         
        local_tmr_voter(481)  <=    (tmr_registers(0)(481) and tmr_registers(1)(481)) or                                                             
                            (tmr_registers(1)(481) and tmr_registers(2)(481)) or                                                             
                            (tmr_registers(0)(481) and tmr_registers(2)(481));                                                               
                                                                                                                                         
        local_tmr_voter(482)  <=    (tmr_registers(0)(482) and tmr_registers(1)(482)) or                                                             
                            (tmr_registers(1)(482) and tmr_registers(2)(482)) or                                                             
                            (tmr_registers(0)(482) and tmr_registers(2)(482));                                                               
                                                                                                                                         
        local_tmr_voter(483)  <=    (tmr_registers(0)(483) and tmr_registers(1)(483)) or                                                             
                            (tmr_registers(1)(483) and tmr_registers(2)(483)) or                                                             
                            (tmr_registers(0)(483) and tmr_registers(2)(483));                                                               
                                                                                                                                         
        local_tmr_voter(484)  <=    (tmr_registers(0)(484) and tmr_registers(1)(484)) or                                                             
                            (tmr_registers(1)(484) and tmr_registers(2)(484)) or                                                             
                            (tmr_registers(0)(484) and tmr_registers(2)(484));                                                               
                                                                                                                                         
        local_tmr_voter(485)  <=    (tmr_registers(0)(485) and tmr_registers(1)(485)) or                                                             
                            (tmr_registers(1)(485) and tmr_registers(2)(485)) or                                                             
                            (tmr_registers(0)(485) and tmr_registers(2)(485));                                                               
                                                                                                                                         
        local_tmr_voter(486)  <=    (tmr_registers(0)(486) and tmr_registers(1)(486)) or                                                             
                            (tmr_registers(1)(486) and tmr_registers(2)(486)) or                                                             
                            (tmr_registers(0)(486) and tmr_registers(2)(486));                                                               
                                                                                                                                         
        local_tmr_voter(487)  <=    (tmr_registers(0)(487) and tmr_registers(1)(487)) or                                                             
                            (tmr_registers(1)(487) and tmr_registers(2)(487)) or                                                             
                            (tmr_registers(0)(487) and tmr_registers(2)(487));                                                               
                                                                                                                                         
        local_tmr_voter(488)  <=    (tmr_registers(0)(488) and tmr_registers(1)(488)) or                                                             
                            (tmr_registers(1)(488) and tmr_registers(2)(488)) or                                                             
                            (tmr_registers(0)(488) and tmr_registers(2)(488));                                                               
                                                                                                                                         
        local_tmr_voter(489)  <=    (tmr_registers(0)(489) and tmr_registers(1)(489)) or                                                             
                            (tmr_registers(1)(489) and tmr_registers(2)(489)) or                                                             
                            (tmr_registers(0)(489) and tmr_registers(2)(489));                                                               
                                                                                                                                         
        local_tmr_voter(490)  <=    (tmr_registers(0)(490) and tmr_registers(1)(490)) or                                                             
                            (tmr_registers(1)(490) and tmr_registers(2)(490)) or                                                             
                            (tmr_registers(0)(490) and tmr_registers(2)(490));                                                               
                                                                                                                                         
        local_tmr_voter(491)  <=    (tmr_registers(0)(491) and tmr_registers(1)(491)) or                                                             
                            (tmr_registers(1)(491) and tmr_registers(2)(491)) or                                                             
                            (tmr_registers(0)(491) and tmr_registers(2)(491));                                                               
                                                                                                                                         
        local_tmr_voter(492)  <=    (tmr_registers(0)(492) and tmr_registers(1)(492)) or                                                             
                            (tmr_registers(1)(492) and tmr_registers(2)(492)) or                                                             
                            (tmr_registers(0)(492) and tmr_registers(2)(492));                                                               
                                                                                                                                         
        local_tmr_voter(493)  <=    (tmr_registers(0)(493) and tmr_registers(1)(493)) or                                                             
                            (tmr_registers(1)(493) and tmr_registers(2)(493)) or                                                             
                            (tmr_registers(0)(493) and tmr_registers(2)(493));                                                               
                                                                                                                                         
        local_tmr_voter(494)  <=    (tmr_registers(0)(494) and tmr_registers(1)(494)) or                                                             
                            (tmr_registers(1)(494) and tmr_registers(2)(494)) or                                                             
                            (tmr_registers(0)(494) and tmr_registers(2)(494));                                                               
                                                                                                                                         
        local_tmr_voter(495)  <=    (tmr_registers(0)(495) and tmr_registers(1)(495)) or                                                             
                            (tmr_registers(1)(495) and tmr_registers(2)(495)) or                                                             
                            (tmr_registers(0)(495) and tmr_registers(2)(495));                                                               
                                                                                                                                         
        local_tmr_voter(496)  <=    (tmr_registers(0)(496) and tmr_registers(1)(496)) or                                                             
                            (tmr_registers(1)(496) and tmr_registers(2)(496)) or                                                             
                            (tmr_registers(0)(496) and tmr_registers(2)(496));                                                               
                                                                                                                                         
        local_tmr_voter(497)  <=    (tmr_registers(0)(497) and tmr_registers(1)(497)) or                                                             
                            (tmr_registers(1)(497) and tmr_registers(2)(497)) or                                                             
                            (tmr_registers(0)(497) and tmr_registers(2)(497));                                                               
                                                                                                                                         
        local_tmr_voter(498)  <=    (tmr_registers(0)(498) and tmr_registers(1)(498)) or                                                             
                            (tmr_registers(1)(498) and tmr_registers(2)(498)) or                                                             
                            (tmr_registers(0)(498) and tmr_registers(2)(498));                                                               
                                                                                                                                         
        local_tmr_voter(499)  <=    (tmr_registers(0)(499) and tmr_registers(1)(499)) or                                                             
                            (tmr_registers(1)(499) and tmr_registers(2)(499)) or                                                             
                            (tmr_registers(0)(499) and tmr_registers(2)(499));                                                               
                                                                                                                                         
        local_tmr_voter(500)  <=    (tmr_registers(0)(500) and tmr_registers(1)(500)) or                                                             
                            (tmr_registers(1)(500) and tmr_registers(2)(500)) or                                                             
                            (tmr_registers(0)(500) and tmr_registers(2)(500));                                                               
                                                                                                                                         
        local_tmr_voter(501)  <=    (tmr_registers(0)(501) and tmr_registers(1)(501)) or                                                             
                            (tmr_registers(1)(501) and tmr_registers(2)(501)) or                                                             
                            (tmr_registers(0)(501) and tmr_registers(2)(501));                                                               
                                                                                                                                         
        local_tmr_voter(502)  <=    (tmr_registers(0)(502) and tmr_registers(1)(502)) or                                                             
                            (tmr_registers(1)(502) and tmr_registers(2)(502)) or                                                             
                            (tmr_registers(0)(502) and tmr_registers(2)(502));                                                               
                                                                                                                                         
        local_tmr_voter(503)  <=    (tmr_registers(0)(503) and tmr_registers(1)(503)) or                                                             
                            (tmr_registers(1)(503) and tmr_registers(2)(503)) or                                                             
                            (tmr_registers(0)(503) and tmr_registers(2)(503));                                                               
                                                                                                                                         
        local_tmr_voter(504)  <=    (tmr_registers(0)(504) and tmr_registers(1)(504)) or                                                             
                            (tmr_registers(1)(504) and tmr_registers(2)(504)) or                                                             
                            (tmr_registers(0)(504) and tmr_registers(2)(504));                                                               
                                                                                                                                         
        local_tmr_voter(505)  <=    (tmr_registers(0)(505) and tmr_registers(1)(505)) or                                                             
                            (tmr_registers(1)(505) and tmr_registers(2)(505)) or                                                             
                            (tmr_registers(0)(505) and tmr_registers(2)(505));                                                               
                                                                                                                                         
        local_tmr_voter(506)  <=    (tmr_registers(0)(506) and tmr_registers(1)(506)) or                                                             
                            (tmr_registers(1)(506) and tmr_registers(2)(506)) or                                                             
                            (tmr_registers(0)(506) and tmr_registers(2)(506));                                                               
                                                                                                                                         
        local_tmr_voter(507)  <=    (tmr_registers(0)(507) and tmr_registers(1)(507)) or                                                             
                            (tmr_registers(1)(507) and tmr_registers(2)(507)) or                                                             
                            (tmr_registers(0)(507) and tmr_registers(2)(507));                                                               
                                                                                                                                         
        local_tmr_voter(508)  <=    (tmr_registers(0)(508) and tmr_registers(1)(508)) or                                                             
                            (tmr_registers(1)(508) and tmr_registers(2)(508)) or                                                             
                            (tmr_registers(0)(508) and tmr_registers(2)(508));                                                               
                                                                                                                                         
        local_tmr_voter(509)  <=    (tmr_registers(0)(509) and tmr_registers(1)(509)) or                                                             
                            (tmr_registers(1)(509) and tmr_registers(2)(509)) or                                                             
                            (tmr_registers(0)(509) and tmr_registers(2)(509));                                                               
                                                                                                                                         
        local_tmr_voter(510)  <=    (tmr_registers(0)(510) and tmr_registers(1)(510)) or                                                             
                            (tmr_registers(1)(510) and tmr_registers(2)(510)) or                                                             
                            (tmr_registers(0)(510) and tmr_registers(2)(510));                                                               
                                                                                                                                         
        local_tmr_voter(511)  <=    (tmr_registers(0)(511) and tmr_registers(1)(511)) or                                                             
                            (tmr_registers(1)(511) and tmr_registers(2)(511)) or                                                             
                            (tmr_registers(0)(511) and tmr_registers(2)(511));                                                               
                                                                                                                                         
        local_tmr_voter(512)  <=    (tmr_registers(0)(512) and tmr_registers(1)(512)) or                                                             
                            (tmr_registers(1)(512) and tmr_registers(2)(512)) or                                                             
                            (tmr_registers(0)(512) and tmr_registers(2)(512));                                                               
                                                                                                                                         
        local_tmr_voter(513)  <=    (tmr_registers(0)(513) and tmr_registers(1)(513)) or                                                             
                            (tmr_registers(1)(513) and tmr_registers(2)(513)) or                                                             
                            (tmr_registers(0)(513) and tmr_registers(2)(513));                                                               
                                                                                                                                         
        local_tmr_voter(514)  <=    (tmr_registers(0)(514) and tmr_registers(1)(514)) or                                                             
                            (tmr_registers(1)(514) and tmr_registers(2)(514)) or                                                             
                            (tmr_registers(0)(514) and tmr_registers(2)(514));                                                               
                                                                                                                                         
        local_tmr_voter(515)  <=    (tmr_registers(0)(515) and tmr_registers(1)(515)) or                                                             
                            (tmr_registers(1)(515) and tmr_registers(2)(515)) or                                                             
                            (tmr_registers(0)(515) and tmr_registers(2)(515));                                                               
                                                                                                                                         
        local_tmr_voter(516)  <=    (tmr_registers(0)(516) and tmr_registers(1)(516)) or                                                             
                            (tmr_registers(1)(516) and tmr_registers(2)(516)) or                                                             
                            (tmr_registers(0)(516) and tmr_registers(2)(516));                                                               
                                                                                                                                         
        local_tmr_voter(517)  <=    (tmr_registers(0)(517) and tmr_registers(1)(517)) or                                                             
                            (tmr_registers(1)(517) and tmr_registers(2)(517)) or                                                             
                            (tmr_registers(0)(517) and tmr_registers(2)(517));                                                               
                                                                                                                                         
        local_tmr_voter(518)  <=    (tmr_registers(0)(518) and tmr_registers(1)(518)) or                                                             
                            (tmr_registers(1)(518) and tmr_registers(2)(518)) or                                                             
                            (tmr_registers(0)(518) and tmr_registers(2)(518));                                                               
                                                                                                                                         
        local_tmr_voter(519)  <=    (tmr_registers(0)(519) and tmr_registers(1)(519)) or                                                             
                            (tmr_registers(1)(519) and tmr_registers(2)(519)) or                                                             
                            (tmr_registers(0)(519) and tmr_registers(2)(519));                                                               
                                                                                                                                         
        local_tmr_voter(520)  <=    (tmr_registers(0)(520) and tmr_registers(1)(520)) or                                                             
                            (tmr_registers(1)(520) and tmr_registers(2)(520)) or                                                             
                            (tmr_registers(0)(520) and tmr_registers(2)(520));                                                               
                                                                                                                                         
        local_tmr_voter(521)  <=    (tmr_registers(0)(521) and tmr_registers(1)(521)) or                                                             
                            (tmr_registers(1)(521) and tmr_registers(2)(521)) or                                                             
                            (tmr_registers(0)(521) and tmr_registers(2)(521));                                                               
                                                                                                                                         
        local_tmr_voter(522)  <=    (tmr_registers(0)(522) and tmr_registers(1)(522)) or                                                             
                            (tmr_registers(1)(522) and tmr_registers(2)(522)) or                                                             
                            (tmr_registers(0)(522) and tmr_registers(2)(522));                                                               
                                                                                                                                         
        local_tmr_voter(523)  <=    (tmr_registers(0)(523) and tmr_registers(1)(523)) or                                                             
                            (tmr_registers(1)(523) and tmr_registers(2)(523)) or                                                             
                            (tmr_registers(0)(523) and tmr_registers(2)(523));                                                               
                                                                                                                                         
        local_tmr_voter(524)  <=    (tmr_registers(0)(524) and tmr_registers(1)(524)) or                                                             
                            (tmr_registers(1)(524) and tmr_registers(2)(524)) or                                                             
                            (tmr_registers(0)(524) and tmr_registers(2)(524));                                                               
                                                                                                                                         
        local_tmr_voter(525)  <=    (tmr_registers(0)(525) and tmr_registers(1)(525)) or                                                             
                            (tmr_registers(1)(525) and tmr_registers(2)(525)) or                                                             
                            (tmr_registers(0)(525) and tmr_registers(2)(525));                                                               
                                                                                                                                         
        local_tmr_voter(526)  <=    (tmr_registers(0)(526) and tmr_registers(1)(526)) or                                                             
                            (tmr_registers(1)(526) and tmr_registers(2)(526)) or                                                             
                            (tmr_registers(0)(526) and tmr_registers(2)(526));                                                               
                                                                                                                                         
        local_tmr_voter(527)  <=    (tmr_registers(0)(527) and tmr_registers(1)(527)) or                                                             
                            (tmr_registers(1)(527) and tmr_registers(2)(527)) or                                                             
                            (tmr_registers(0)(527) and tmr_registers(2)(527));                                                               
                                                                                                                                         
        local_tmr_voter(528)  <=    (tmr_registers(0)(528) and tmr_registers(1)(528)) or                                                             
                            (tmr_registers(1)(528) and tmr_registers(2)(528)) or                                                             
                            (tmr_registers(0)(528) and tmr_registers(2)(528));                                                               
                                                                                                                                         
        local_tmr_voter(529)  <=    (tmr_registers(0)(529) and tmr_registers(1)(529)) or                                                             
                            (tmr_registers(1)(529) and tmr_registers(2)(529)) or                                                             
                            (tmr_registers(0)(529) and tmr_registers(2)(529));                                                               
                                                                                                                                         
        local_tmr_voter(530)  <=    (tmr_registers(0)(530) and tmr_registers(1)(530)) or                                                             
                            (tmr_registers(1)(530) and tmr_registers(2)(530)) or                                                             
                            (tmr_registers(0)(530) and tmr_registers(2)(530));                                                               
                                                                                                                                         
        local_tmr_voter(531)  <=    (tmr_registers(0)(531) and tmr_registers(1)(531)) or                                                             
                            (tmr_registers(1)(531) and tmr_registers(2)(531)) or                                                             
                            (tmr_registers(0)(531) and tmr_registers(2)(531));                                                               
                                                                                                                                         
        local_tmr_voter(532)  <=    (tmr_registers(0)(532) and tmr_registers(1)(532)) or                                                             
                            (tmr_registers(1)(532) and tmr_registers(2)(532)) or                                                             
                            (tmr_registers(0)(532) and tmr_registers(2)(532));                                                               
                                                                                                                                         
        local_tmr_voter(533)  <=    (tmr_registers(0)(533) and tmr_registers(1)(533)) or                                                             
                            (tmr_registers(1)(533) and tmr_registers(2)(533)) or                                                             
                            (tmr_registers(0)(533) and tmr_registers(2)(533));                                                               
                                                                                                                                         
        local_tmr_voter(534)  <=    (tmr_registers(0)(534) and tmr_registers(1)(534)) or                                                             
                            (tmr_registers(1)(534) and tmr_registers(2)(534)) or                                                             
                            (tmr_registers(0)(534) and tmr_registers(2)(534));                                                               
                                                                                                                                         
        local_tmr_voter(535)  <=    (tmr_registers(0)(535) and tmr_registers(1)(535)) or                                                             
                            (tmr_registers(1)(535) and tmr_registers(2)(535)) or                                                             
                            (tmr_registers(0)(535) and tmr_registers(2)(535));                                                               
                                                                                                                                         
        local_tmr_voter(536)  <=    (tmr_registers(0)(536) and tmr_registers(1)(536)) or                                                             
                            (tmr_registers(1)(536) and tmr_registers(2)(536)) or                                                             
                            (tmr_registers(0)(536) and tmr_registers(2)(536));                                                               
                                                                                                                                         
        local_tmr_voter(537)  <=    (tmr_registers(0)(537) and tmr_registers(1)(537)) or                                                             
                            (tmr_registers(1)(537) and tmr_registers(2)(537)) or                                                             
                            (tmr_registers(0)(537) and tmr_registers(2)(537));                                                               
                                                                                                                                         
        local_tmr_voter(538)  <=    (tmr_registers(0)(538) and tmr_registers(1)(538)) or                                                             
                            (tmr_registers(1)(538) and tmr_registers(2)(538)) or                                                             
                            (tmr_registers(0)(538) and tmr_registers(2)(538));                                                               
                                                                                                                                         
        local_tmr_voter(539)  <=    (tmr_registers(0)(539) and tmr_registers(1)(539)) or                                                             
                            (tmr_registers(1)(539) and tmr_registers(2)(539)) or                                                             
                            (tmr_registers(0)(539) and tmr_registers(2)(539));                                                               
                                                                                                                                         
        local_tmr_voter(540)  <=    (tmr_registers(0)(540) and tmr_registers(1)(540)) or                                                             
                            (tmr_registers(1)(540) and tmr_registers(2)(540)) or                                                             
                            (tmr_registers(0)(540) and tmr_registers(2)(540));                                                               
                                                                                                                                         
        local_tmr_voter(541)  <=    (tmr_registers(0)(541) and tmr_registers(1)(541)) or                                                             
                            (tmr_registers(1)(541) and tmr_registers(2)(541)) or                                                             
                            (tmr_registers(0)(541) and tmr_registers(2)(541));                                                               
                                                                                                                                         
        local_tmr_voter(542)  <=    (tmr_registers(0)(542) and tmr_registers(1)(542)) or                                                             
                            (tmr_registers(1)(542) and tmr_registers(2)(542)) or                                                             
                            (tmr_registers(0)(542) and tmr_registers(2)(542));                                                               
                                                                                                                                         
        local_tmr_voter(543)  <=    (tmr_registers(0)(543) and tmr_registers(1)(543)) or                                                             
                            (tmr_registers(1)(543) and tmr_registers(2)(543)) or                                                             
                            (tmr_registers(0)(543) and tmr_registers(2)(543));                                                               
                                                                                                                                         
        local_tmr_voter(544)  <=    (tmr_registers(0)(544) and tmr_registers(1)(544)) or                                                             
                            (tmr_registers(1)(544) and tmr_registers(2)(544)) or                                                             
                            (tmr_registers(0)(544) and tmr_registers(2)(544));                                                               
                                                                                                                                         
        local_tmr_voter(545)  <=    (tmr_registers(0)(545) and tmr_registers(1)(545)) or                                                             
                            (tmr_registers(1)(545) and tmr_registers(2)(545)) or                                                             
                            (tmr_registers(0)(545) and tmr_registers(2)(545));                                                               
                                                                                                                                         
        local_tmr_voter(546)  <=    (tmr_registers(0)(546) and tmr_registers(1)(546)) or                                                             
                            (tmr_registers(1)(546) and tmr_registers(2)(546)) or                                                             
                            (tmr_registers(0)(546) and tmr_registers(2)(546));                                                               
                                                                                                                                         
        local_tmr_voter(547)  <=    (tmr_registers(0)(547) and tmr_registers(1)(547)) or                                                             
                            (tmr_registers(1)(547) and tmr_registers(2)(547)) or                                                             
                            (tmr_registers(0)(547) and tmr_registers(2)(547));                                                               
                                                                                                                                         
        local_tmr_voter(548)  <=    (tmr_registers(0)(548) and tmr_registers(1)(548)) or                                                             
                            (tmr_registers(1)(548) and tmr_registers(2)(548)) or                                                             
                            (tmr_registers(0)(548) and tmr_registers(2)(548));                                                               
                                                                                                                                         
        local_tmr_voter(549)  <=    (tmr_registers(0)(549) and tmr_registers(1)(549)) or                                                             
                            (tmr_registers(1)(549) and tmr_registers(2)(549)) or                                                             
                            (tmr_registers(0)(549) and tmr_registers(2)(549));                                                               
                                                                                                                                         
        local_tmr_voter(550)  <=    (tmr_registers(0)(550) and tmr_registers(1)(550)) or                                                             
                            (tmr_registers(1)(550) and tmr_registers(2)(550)) or                                                             
                            (tmr_registers(0)(550) and tmr_registers(2)(550));                                                               
                                                                                                                                         
        local_tmr_voter(551)  <=    (tmr_registers(0)(551) and tmr_registers(1)(551)) or                                                             
                            (tmr_registers(1)(551) and tmr_registers(2)(551)) or                                                             
                            (tmr_registers(0)(551) and tmr_registers(2)(551));                                                               
                                                                                                                                         
        local_tmr_voter(552)  <=    (tmr_registers(0)(552) and tmr_registers(1)(552)) or                                                             
                            (tmr_registers(1)(552) and tmr_registers(2)(552)) or                                                             
                            (tmr_registers(0)(552) and tmr_registers(2)(552));                                                               
                                                                                                                                         
        local_tmr_voter(553)  <=    (tmr_registers(0)(553) and tmr_registers(1)(553)) or                                                             
                            (tmr_registers(1)(553) and tmr_registers(2)(553)) or                                                             
                            (tmr_registers(0)(553) and tmr_registers(2)(553));                                                               
                                                                                                                                         
        local_tmr_voter(554)  <=    (tmr_registers(0)(554) and tmr_registers(1)(554)) or                                                             
                            (tmr_registers(1)(554) and tmr_registers(2)(554)) or                                                             
                            (tmr_registers(0)(554) and tmr_registers(2)(554));                                                               
                                                                                                                                         
        local_tmr_voter(555)  <=    (tmr_registers(0)(555) and tmr_registers(1)(555)) or                                                             
                            (tmr_registers(1)(555) and tmr_registers(2)(555)) or                                                             
                            (tmr_registers(0)(555) and tmr_registers(2)(555));                                                               
                                                                                                                                         
        local_tmr_voter(556)  <=    (tmr_registers(0)(556) and tmr_registers(1)(556)) or                                                             
                            (tmr_registers(1)(556) and tmr_registers(2)(556)) or                                                             
                            (tmr_registers(0)(556) and tmr_registers(2)(556));                                                               
                                                                                                                                         
        local_tmr_voter(557)  <=    (tmr_registers(0)(557) and tmr_registers(1)(557)) or                                                             
                            (tmr_registers(1)(557) and tmr_registers(2)(557)) or                                                             
                            (tmr_registers(0)(557) and tmr_registers(2)(557));                                                               
                                                                                                                                         
        local_tmr_voter(558)  <=    (tmr_registers(0)(558) and tmr_registers(1)(558)) or                                                             
                            (tmr_registers(1)(558) and tmr_registers(2)(558)) or                                                             
                            (tmr_registers(0)(558) and tmr_registers(2)(558));                                                               
                                                                                                                                         
        local_tmr_voter(559)  <=    (tmr_registers(0)(559) and tmr_registers(1)(559)) or                                                             
                            (tmr_registers(1)(559) and tmr_registers(2)(559)) or                                                             
                            (tmr_registers(0)(559) and tmr_registers(2)(559));                                                               
                                                                                                                                         
        local_tmr_voter(560)  <=    (tmr_registers(0)(560) and tmr_registers(1)(560)) or                                                             
                            (tmr_registers(1)(560) and tmr_registers(2)(560)) or                                                             
                            (tmr_registers(0)(560) and tmr_registers(2)(560));                                                               
                                                                                                                                         
        local_tmr_voter(561)  <=    (tmr_registers(0)(561) and tmr_registers(1)(561)) or                                                             
                            (tmr_registers(1)(561) and tmr_registers(2)(561)) or                                                             
                            (tmr_registers(0)(561) and tmr_registers(2)(561));                                                               
                                                                                                                                         
        local_tmr_voter(562)  <=    (tmr_registers(0)(562) and tmr_registers(1)(562)) or                                                             
                            (tmr_registers(1)(562) and tmr_registers(2)(562)) or                                                             
                            (tmr_registers(0)(562) and tmr_registers(2)(562));                                                               
                                                                                                                                         
        local_tmr_voter(563)  <=    (tmr_registers(0)(563) and tmr_registers(1)(563)) or                                                             
                            (tmr_registers(1)(563) and tmr_registers(2)(563)) or                                                             
                            (tmr_registers(0)(563) and tmr_registers(2)(563));                                                               
                                                                                                                                         
        local_tmr_voter(564)  <=    (tmr_registers(0)(564) and tmr_registers(1)(564)) or                                                             
                            (tmr_registers(1)(564) and tmr_registers(2)(564)) or                                                             
                            (tmr_registers(0)(564) and tmr_registers(2)(564));                                                               
                                                                                                                                         
        local_tmr_voter(565)  <=    (tmr_registers(0)(565) and tmr_registers(1)(565)) or                                                             
                            (tmr_registers(1)(565) and tmr_registers(2)(565)) or                                                             
                            (tmr_registers(0)(565) and tmr_registers(2)(565));                                                               
                                                                                                                                         
        local_tmr_voter(566)  <=    (tmr_registers(0)(566) and tmr_registers(1)(566)) or                                                             
                            (tmr_registers(1)(566) and tmr_registers(2)(566)) or                                                             
                            (tmr_registers(0)(566) and tmr_registers(2)(566));                                                               
                                                                                                                                         
        local_tmr_voter(567)  <=    (tmr_registers(0)(567) and tmr_registers(1)(567)) or                                                             
                            (tmr_registers(1)(567) and tmr_registers(2)(567)) or                                                             
                            (tmr_registers(0)(567) and tmr_registers(2)(567));                                                               
                                                                                                                                         
        local_tmr_voter(568)  <=    (tmr_registers(0)(568) and tmr_registers(1)(568)) or                                                             
                            (tmr_registers(1)(568) and tmr_registers(2)(568)) or                                                             
                            (tmr_registers(0)(568) and tmr_registers(2)(568));                                                               
                                                                                                                                         
        local_tmr_voter(569)  <=    (tmr_registers(0)(569) and tmr_registers(1)(569)) or                                                             
                            (tmr_registers(1)(569) and tmr_registers(2)(569)) or                                                             
                            (tmr_registers(0)(569) and tmr_registers(2)(569));                                                               
                                                                                                                                         
        local_tmr_voter(570)  <=    (tmr_registers(0)(570) and tmr_registers(1)(570)) or                                                             
                            (tmr_registers(1)(570) and tmr_registers(2)(570)) or                                                             
                            (tmr_registers(0)(570) and tmr_registers(2)(570));                                                               
                                                                                                                                         
        local_tmr_voter(571)  <=    (tmr_registers(0)(571) and tmr_registers(1)(571)) or                                                             
                            (tmr_registers(1)(571) and tmr_registers(2)(571)) or                                                             
                            (tmr_registers(0)(571) and tmr_registers(2)(571));                                                               
                                                                                                                                         
        local_tmr_voter(572)  <=    (tmr_registers(0)(572) and tmr_registers(1)(572)) or                                                             
                            (tmr_registers(1)(572) and tmr_registers(2)(572)) or                                                             
                            (tmr_registers(0)(572) and tmr_registers(2)(572));                                                               
                                                                                                                                         
        local_tmr_voter(573)  <=    (tmr_registers(0)(573) and tmr_registers(1)(573)) or                                                             
                            (tmr_registers(1)(573) and tmr_registers(2)(573)) or                                                             
                            (tmr_registers(0)(573) and tmr_registers(2)(573));                                                               
                                                                                                                                         
        local_tmr_voter(574)  <=    (tmr_registers(0)(574) and tmr_registers(1)(574)) or                                                             
                            (tmr_registers(1)(574) and tmr_registers(2)(574)) or                                                             
                            (tmr_registers(0)(574) and tmr_registers(2)(574));                                                               
                                                                                                                                         
        local_tmr_voter(575)  <=    (tmr_registers(0)(575) and tmr_registers(1)(575)) or                                                             
                            (tmr_registers(1)(575) and tmr_registers(2)(575)) or                                                             
                            (tmr_registers(0)(575) and tmr_registers(2)(575));                                                               
                                                                                                                                         
        local_tmr_voter(576)  <=    (tmr_registers(0)(576) and tmr_registers(1)(576)) or                                                             
                            (tmr_registers(1)(576) and tmr_registers(2)(576)) or                                                             
                            (tmr_registers(0)(576) and tmr_registers(2)(576));                                                               
                                                                                                                                         
        local_tmr_voter(577)  <=    (tmr_registers(0)(577) and tmr_registers(1)(577)) or                                                             
                            (tmr_registers(1)(577) and tmr_registers(2)(577)) or                                                             
                            (tmr_registers(0)(577) and tmr_registers(2)(577));                                                               
                                                                                                                                         
        local_tmr_voter(578)  <=    (tmr_registers(0)(578) and tmr_registers(1)(578)) or                                                             
                            (tmr_registers(1)(578) and tmr_registers(2)(578)) or                                                             
                            (tmr_registers(0)(578) and tmr_registers(2)(578));                                                               
                                                                                                                                         
        local_tmr_voter(579)  <=    (tmr_registers(0)(579) and tmr_registers(1)(579)) or                                                             
                            (tmr_registers(1)(579) and tmr_registers(2)(579)) or                                                             
                            (tmr_registers(0)(579) and tmr_registers(2)(579));                                                               
                                                                                                                                         
        local_tmr_voter(580)  <=    (tmr_registers(0)(580) and tmr_registers(1)(580)) or                                                             
                            (tmr_registers(1)(580) and tmr_registers(2)(580)) or                                                             
                            (tmr_registers(0)(580) and tmr_registers(2)(580));                                                               
                                                                                                                                         
        local_tmr_voter(581)  <=    (tmr_registers(0)(581) and tmr_registers(1)(581)) or                                                             
                            (tmr_registers(1)(581) and tmr_registers(2)(581)) or                                                             
                            (tmr_registers(0)(581) and tmr_registers(2)(581));                                                               
                                                                                                                                         
        local_tmr_voter(582)  <=    (tmr_registers(0)(582) and tmr_registers(1)(582)) or                                                             
                            (tmr_registers(1)(582) and tmr_registers(2)(582)) or                                                             
                            (tmr_registers(0)(582) and tmr_registers(2)(582));                                                               
                                                                                                                                         
        local_tmr_voter(583)  <=    (tmr_registers(0)(583) and tmr_registers(1)(583)) or                                                             
                            (tmr_registers(1)(583) and tmr_registers(2)(583)) or                                                             
                            (tmr_registers(0)(583) and tmr_registers(2)(583));                                                               
                                                                                                                                         
        local_tmr_voter(584)  <=    (tmr_registers(0)(584) and tmr_registers(1)(584)) or                                                             
                            (tmr_registers(1)(584) and tmr_registers(2)(584)) or                                                             
                            (tmr_registers(0)(584) and tmr_registers(2)(584));                                                               
                                                                                                                                         
        local_tmr_voter(585)  <=    (tmr_registers(0)(585) and tmr_registers(1)(585)) or                                                             
                            (tmr_registers(1)(585) and tmr_registers(2)(585)) or                                                             
                            (tmr_registers(0)(585) and tmr_registers(2)(585));                                                               
                                                                                                                                         
        local_tmr_voter(586)  <=    (tmr_registers(0)(586) and tmr_registers(1)(586)) or                                                             
                            (tmr_registers(1)(586) and tmr_registers(2)(586)) or                                                             
                            (tmr_registers(0)(586) and tmr_registers(2)(586));                                                               
                                                                                                                                         
        local_tmr_voter(587)  <=    (tmr_registers(0)(587) and tmr_registers(1)(587)) or                                                             
                            (tmr_registers(1)(587) and tmr_registers(2)(587)) or                                                             
                            (tmr_registers(0)(587) and tmr_registers(2)(587));                                                               
                                                                                                                                         
        local_tmr_voter(588)  <=    (tmr_registers(0)(588) and tmr_registers(1)(588)) or                                                             
                            (tmr_registers(1)(588) and tmr_registers(2)(588)) or                                                             
                            (tmr_registers(0)(588) and tmr_registers(2)(588));                                                               
                                                                                                                                         
        local_tmr_voter(589)  <=    (tmr_registers(0)(589) and tmr_registers(1)(589)) or                                                             
                            (tmr_registers(1)(589) and tmr_registers(2)(589)) or                                                             
                            (tmr_registers(0)(589) and tmr_registers(2)(589));                                                               
                                                                                                                                         
        local_tmr_voter(590)  <=    (tmr_registers(0)(590) and tmr_registers(1)(590)) or                                                             
                            (tmr_registers(1)(590) and tmr_registers(2)(590)) or                                                             
                            (tmr_registers(0)(590) and tmr_registers(2)(590));                                                               
                                                                                                                                         
        local_tmr_voter(591)  <=    (tmr_registers(0)(591) and tmr_registers(1)(591)) or                                                             
                            (tmr_registers(1)(591) and tmr_registers(2)(591)) or                                                             
                            (tmr_registers(0)(591) and tmr_registers(2)(591));                                                               
                                                                                                                                         
        local_tmr_voter(592)  <=    (tmr_registers(0)(592) and tmr_registers(1)(592)) or                                                             
                            (tmr_registers(1)(592) and tmr_registers(2)(592)) or                                                             
                            (tmr_registers(0)(592) and tmr_registers(2)(592));                                                               
                                                                                                                                         
        local_tmr_voter(593)  <=    (tmr_registers(0)(593) and tmr_registers(1)(593)) or                                                             
                            (tmr_registers(1)(593) and tmr_registers(2)(593)) or                                                             
                            (tmr_registers(0)(593) and tmr_registers(2)(593));                                                               
                                                                                                                                         
        local_tmr_voter(594)  <=    (tmr_registers(0)(594) and tmr_registers(1)(594)) or                                                             
                            (tmr_registers(1)(594) and tmr_registers(2)(594)) or                                                             
                            (tmr_registers(0)(594) and tmr_registers(2)(594));                                                               
                                                                                                                                         
        local_tmr_voter(595)  <=    (tmr_registers(0)(595) and tmr_registers(1)(595)) or                                                             
                            (tmr_registers(1)(595) and tmr_registers(2)(595)) or                                                             
                            (tmr_registers(0)(595) and tmr_registers(2)(595));                                                               
                                                                                                                                         
        local_tmr_voter(596)  <=    (tmr_registers(0)(596) and tmr_registers(1)(596)) or                                                             
                            (tmr_registers(1)(596) and tmr_registers(2)(596)) or                                                             
                            (tmr_registers(0)(596) and tmr_registers(2)(596));                                                               
                                                                                                                                         
        local_tmr_voter(597)  <=    (tmr_registers(0)(597) and tmr_registers(1)(597)) or                                                             
                            (tmr_registers(1)(597) and tmr_registers(2)(597)) or                                                             
                            (tmr_registers(0)(597) and tmr_registers(2)(597));                                                               
                                                                                                                                         
        local_tmr_voter(598)  <=    (tmr_registers(0)(598) and tmr_registers(1)(598)) or                                                             
                            (tmr_registers(1)(598) and tmr_registers(2)(598)) or                                                             
                            (tmr_registers(0)(598) and tmr_registers(2)(598));                                                               
                                                                                                                                         
        local_tmr_voter(599)  <=    (tmr_registers(0)(599) and tmr_registers(1)(599)) or                                                             
                            (tmr_registers(1)(599) and tmr_registers(2)(599)) or                                                             
                            (tmr_registers(0)(599) and tmr_registers(2)(599));                                                               
                                                                                                                                         
        local_tmr_voter(600)  <=    (tmr_registers(0)(600) and tmr_registers(1)(600)) or                                                             
                            (tmr_registers(1)(600) and tmr_registers(2)(600)) or                                                             
                            (tmr_registers(0)(600) and tmr_registers(2)(600));                                                               
                                                                                                                                         
        local_tmr_voter(601)  <=    (tmr_registers(0)(601) and tmr_registers(1)(601)) or                                                             
                            (tmr_registers(1)(601) and tmr_registers(2)(601)) or                                                             
                            (tmr_registers(0)(601) and tmr_registers(2)(601));                                                               
                                                                                                                                         
        local_tmr_voter(602)  <=    (tmr_registers(0)(602) and tmr_registers(1)(602)) or                                                             
                            (tmr_registers(1)(602) and tmr_registers(2)(602)) or                                                             
                            (tmr_registers(0)(602) and tmr_registers(2)(602));                                                               
                                                                                                                                         
        local_tmr_voter(603)  <=    (tmr_registers(0)(603) and tmr_registers(1)(603)) or                                                             
                            (tmr_registers(1)(603) and tmr_registers(2)(603)) or                                                             
                            (tmr_registers(0)(603) and tmr_registers(2)(603));                                                               
                                                                                                                                         
        local_tmr_voter(604)  <=    (tmr_registers(0)(604) and tmr_registers(1)(604)) or                                                             
                            (tmr_registers(1)(604) and tmr_registers(2)(604)) or                                                             
                            (tmr_registers(0)(604) and tmr_registers(2)(604));                                                               
                                                                                                                                         
        local_tmr_voter(605)  <=    (tmr_registers(0)(605) and tmr_registers(1)(605)) or                                                             
                            (tmr_registers(1)(605) and tmr_registers(2)(605)) or                                                             
                            (tmr_registers(0)(605) and tmr_registers(2)(605));                                                               
                                                                                                                                         
        local_tmr_voter(606)  <=    (tmr_registers(0)(606) and tmr_registers(1)(606)) or                                                             
                            (tmr_registers(1)(606) and tmr_registers(2)(606)) or                                                             
                            (tmr_registers(0)(606) and tmr_registers(2)(606));                                                               
                                                                                                                                         
        local_tmr_voter(607)  <=    (tmr_registers(0)(607) and tmr_registers(1)(607)) or                                                             
                            (tmr_registers(1)(607) and tmr_registers(2)(607)) or                                                             
                            (tmr_registers(0)(607) and tmr_registers(2)(607));                                                               
                                                                                                                                         
        local_tmr_voter(608)  <=    (tmr_registers(0)(608) and tmr_registers(1)(608)) or                                                             
                            (tmr_registers(1)(608) and tmr_registers(2)(608)) or                                                             
                            (tmr_registers(0)(608) and tmr_registers(2)(608));                                                               
                                                                                                                                         
        local_tmr_voter(609)  <=    (tmr_registers(0)(609) and tmr_registers(1)(609)) or                                                             
                            (tmr_registers(1)(609) and tmr_registers(2)(609)) or                                                             
                            (tmr_registers(0)(609) and tmr_registers(2)(609));                                                               
                                                                                                                                         
        local_tmr_voter(610)  <=    (tmr_registers(0)(610) and tmr_registers(1)(610)) or                                                             
                            (tmr_registers(1)(610) and tmr_registers(2)(610)) or                                                             
                            (tmr_registers(0)(610) and tmr_registers(2)(610));                                                               
                                                                                                                                         
        local_tmr_voter(611)  <=    (tmr_registers(0)(611) and tmr_registers(1)(611)) or                                                             
                            (tmr_registers(1)(611) and tmr_registers(2)(611)) or                                                             
                            (tmr_registers(0)(611) and tmr_registers(2)(611));                                                               
                                                                                                                                         
        local_tmr_voter(612)  <=    (tmr_registers(0)(612) and tmr_registers(1)(612)) or                                                             
                            (tmr_registers(1)(612) and tmr_registers(2)(612)) or                                                             
                            (tmr_registers(0)(612) and tmr_registers(2)(612));                                                               
                                                                                                                                         
        local_tmr_voter(613)  <=    (tmr_registers(0)(613) and tmr_registers(1)(613)) or                                                             
                            (tmr_registers(1)(613) and tmr_registers(2)(613)) or                                                             
                            (tmr_registers(0)(613) and tmr_registers(2)(613));                                                               
                                                                                                                                         
        local_tmr_voter(614)  <=    (tmr_registers(0)(614) and tmr_registers(1)(614)) or                                                             
                            (tmr_registers(1)(614) and tmr_registers(2)(614)) or                                                             
                            (tmr_registers(0)(614) and tmr_registers(2)(614));                                                               
                                                                                                                                         
        local_tmr_voter(615)  <=    (tmr_registers(0)(615) and tmr_registers(1)(615)) or                                                             
                            (tmr_registers(1)(615) and tmr_registers(2)(615)) or                                                             
                            (tmr_registers(0)(615) and tmr_registers(2)(615));                                                               
                                                                                                                                         
        local_tmr_voter(616)  <=    (tmr_registers(0)(616) and tmr_registers(1)(616)) or                                                             
                            (tmr_registers(1)(616) and tmr_registers(2)(616)) or                                                             
                            (tmr_registers(0)(616) and tmr_registers(2)(616));                                                               
                                                                                                                                         
        local_tmr_voter(617)  <=    (tmr_registers(0)(617) and tmr_registers(1)(617)) or                                                             
                            (tmr_registers(1)(617) and tmr_registers(2)(617)) or                                                             
                            (tmr_registers(0)(617) and tmr_registers(2)(617));                                                               
                                                                                                                                         
        local_tmr_voter(618)  <=    (tmr_registers(0)(618) and tmr_registers(1)(618)) or                                                             
                            (tmr_registers(1)(618) and tmr_registers(2)(618)) or                                                             
                            (tmr_registers(0)(618) and tmr_registers(2)(618));                                                               
                                                                                                                                         
        local_tmr_voter(619)  <=    (tmr_registers(0)(619) and tmr_registers(1)(619)) or                                                             
                            (tmr_registers(1)(619) and tmr_registers(2)(619)) or                                                             
                            (tmr_registers(0)(619) and tmr_registers(2)(619));                                                               
                                                                                                                                         
        local_tmr_voter(620)  <=    (tmr_registers(0)(620) and tmr_registers(1)(620)) or                                                             
                            (tmr_registers(1)(620) and tmr_registers(2)(620)) or                                                             
                            (tmr_registers(0)(620) and tmr_registers(2)(620));                                                               
                                                                                                                                         
        local_tmr_voter(621)  <=    (tmr_registers(0)(621) and tmr_registers(1)(621)) or                                                             
                            (tmr_registers(1)(621) and tmr_registers(2)(621)) or                                                             
                            (tmr_registers(0)(621) and tmr_registers(2)(621));                                                               
                                                                                                                                         
        local_tmr_voter(622)  <=    (tmr_registers(0)(622) and tmr_registers(1)(622)) or                                                             
                            (tmr_registers(1)(622) and tmr_registers(2)(622)) or                                                             
                            (tmr_registers(0)(622) and tmr_registers(2)(622));                                                               
                                                                                                                                         
        local_tmr_voter(623)  <=    (tmr_registers(0)(623) and tmr_registers(1)(623)) or                                                             
                            (tmr_registers(1)(623) and tmr_registers(2)(623)) or                                                             
                            (tmr_registers(0)(623) and tmr_registers(2)(623));                                                               
                                                                                                                                         
        local_tmr_voter(624)  <=    (tmr_registers(0)(624) and tmr_registers(1)(624)) or                                                             
                            (tmr_registers(1)(624) and tmr_registers(2)(624)) or                                                             
                            (tmr_registers(0)(624) and tmr_registers(2)(624));                                                               
                                                                                                                                         
        local_tmr_voter(625)  <=    (tmr_registers(0)(625) and tmr_registers(1)(625)) or                                                             
                            (tmr_registers(1)(625) and tmr_registers(2)(625)) or                                                             
                            (tmr_registers(0)(625) and tmr_registers(2)(625));                                                               
                                                                                                                                         
        local_tmr_voter(626)  <=    (tmr_registers(0)(626) and tmr_registers(1)(626)) or                                                             
                            (tmr_registers(1)(626) and tmr_registers(2)(626)) or                                                             
                            (tmr_registers(0)(626) and tmr_registers(2)(626));                                                               
                                                                                                                                         
        local_tmr_voter(627)  <=    (tmr_registers(0)(627) and tmr_registers(1)(627)) or                                                             
                            (tmr_registers(1)(627) and tmr_registers(2)(627)) or                                                             
                            (tmr_registers(0)(627) and tmr_registers(2)(627));                                                               
                                                                                                                                         
        local_tmr_voter(628)  <=    (tmr_registers(0)(628) and tmr_registers(1)(628)) or                                                             
                            (tmr_registers(1)(628) and tmr_registers(2)(628)) or                                                             
                            (tmr_registers(0)(628) and tmr_registers(2)(628));                                                               
                                                                                                                                         
        local_tmr_voter(629)  <=    (tmr_registers(0)(629) and tmr_registers(1)(629)) or                                                             
                            (tmr_registers(1)(629) and tmr_registers(2)(629)) or                                                             
                            (tmr_registers(0)(629) and tmr_registers(2)(629));                                                               
                                                                                                                                         
        local_tmr_voter(630)  <=    (tmr_registers(0)(630) and tmr_registers(1)(630)) or                                                             
                            (tmr_registers(1)(630) and tmr_registers(2)(630)) or                                                             
                            (tmr_registers(0)(630) and tmr_registers(2)(630));                                                               
                                                                                                                                         
        local_tmr_voter(631)  <=    (tmr_registers(0)(631) and tmr_registers(1)(631)) or                                                             
                            (tmr_registers(1)(631) and tmr_registers(2)(631)) or                                                             
                            (tmr_registers(0)(631) and tmr_registers(2)(631));                                                               
                                                                                                                                         
        local_tmr_voter(632)  <=    (tmr_registers(0)(632) and tmr_registers(1)(632)) or                                                             
                            (tmr_registers(1)(632) and tmr_registers(2)(632)) or                                                             
                            (tmr_registers(0)(632) and tmr_registers(2)(632));                                                               
                                                                                                                                         
        local_tmr_voter(633)  <=    (tmr_registers(0)(633) and tmr_registers(1)(633)) or                                                             
                            (tmr_registers(1)(633) and tmr_registers(2)(633)) or                                                             
                            (tmr_registers(0)(633) and tmr_registers(2)(633));                                                               
                                                                                                                                         
        local_tmr_voter(634)  <=    (tmr_registers(0)(634) and tmr_registers(1)(634)) or                                                             
                            (tmr_registers(1)(634) and tmr_registers(2)(634)) or                                                             
                            (tmr_registers(0)(634) and tmr_registers(2)(634));                                                               
                                                                                                                                         
        local_tmr_voter(635)  <=    (tmr_registers(0)(635) and tmr_registers(1)(635)) or                                                             
                            (tmr_registers(1)(635) and tmr_registers(2)(635)) or                                                             
                            (tmr_registers(0)(635) and tmr_registers(2)(635));                                                               
                                                                                                                                         
        local_tmr_voter(636)  <=    (tmr_registers(0)(636) and tmr_registers(1)(636)) or                                                             
                            (tmr_registers(1)(636) and tmr_registers(2)(636)) or                                                             
                            (tmr_registers(0)(636) and tmr_registers(2)(636));                                                               
                                                                                                                                         
        local_tmr_voter(637)  <=    (tmr_registers(0)(637) and tmr_registers(1)(637)) or                                                             
                            (tmr_registers(1)(637) and tmr_registers(2)(637)) or                                                             
                            (tmr_registers(0)(637) and tmr_registers(2)(637));                                                               
                                                                                                                                         
        local_tmr_voter(638)  <=    (tmr_registers(0)(638) and tmr_registers(1)(638)) or                                                             
                            (tmr_registers(1)(638) and tmr_registers(2)(638)) or                                                             
                            (tmr_registers(0)(638) and tmr_registers(2)(638));                                                               
                                                                                                                                         
        local_tmr_voter(639)  <=    (tmr_registers(0)(639) and tmr_registers(1)(639)) or                                                             
                            (tmr_registers(1)(639) and tmr_registers(2)(639)) or                                                             
                            (tmr_registers(0)(639) and tmr_registers(2)(639));                                                               
                                                                                                                                         
        local_tmr_voter(640)  <=    (tmr_registers(0)(640) and tmr_registers(1)(640)) or                                                             
                            (tmr_registers(1)(640) and tmr_registers(2)(640)) or                                                             
                            (tmr_registers(0)(640) and tmr_registers(2)(640));                                                               
                                                                                                                                         
        local_tmr_voter(641)  <=    (tmr_registers(0)(641) and tmr_registers(1)(641)) or                                                             
                            (tmr_registers(1)(641) and tmr_registers(2)(641)) or                                                             
                            (tmr_registers(0)(641) and tmr_registers(2)(641));                                                               
                                                                                                                                         
        local_tmr_voter(642)  <=    (tmr_registers(0)(642) and tmr_registers(1)(642)) or                                                             
                            (tmr_registers(1)(642) and tmr_registers(2)(642)) or                                                             
                            (tmr_registers(0)(642) and tmr_registers(2)(642));                                                               
                                                                                                                                         
        local_tmr_voter(643)  <=    (tmr_registers(0)(643) and tmr_registers(1)(643)) or                                                             
                            (tmr_registers(1)(643) and tmr_registers(2)(643)) or                                                             
                            (tmr_registers(0)(643) and tmr_registers(2)(643));                                                               
                                                                                                                                         
        local_tmr_voter(644)  <=    (tmr_registers(0)(644) and tmr_registers(1)(644)) or                                                             
                            (tmr_registers(1)(644) and tmr_registers(2)(644)) or                                                             
                            (tmr_registers(0)(644) and tmr_registers(2)(644));                                                               
                                                                                                                                         
        local_tmr_voter(645)  <=    (tmr_registers(0)(645) and tmr_registers(1)(645)) or                                                             
                            (tmr_registers(1)(645) and tmr_registers(2)(645)) or                                                             
                            (tmr_registers(0)(645) and tmr_registers(2)(645));                                                               
                                                                                                                                         
        local_tmr_voter(646)  <=    (tmr_registers(0)(646) and tmr_registers(1)(646)) or                                                             
                            (tmr_registers(1)(646) and tmr_registers(2)(646)) or                                                             
                            (tmr_registers(0)(646) and tmr_registers(2)(646));                                                               
                                                                                                                                         
        local_tmr_voter(647)  <=    (tmr_registers(0)(647) and tmr_registers(1)(647)) or                                                             
                            (tmr_registers(1)(647) and tmr_registers(2)(647)) or                                                             
                            (tmr_registers(0)(647) and tmr_registers(2)(647));                                                               
                                                                                                                                         
        local_tmr_voter(648)  <=    (tmr_registers(0)(648) and tmr_registers(1)(648)) or                                                             
                            (tmr_registers(1)(648) and tmr_registers(2)(648)) or                                                             
                            (tmr_registers(0)(648) and tmr_registers(2)(648));                                                               
                                                                                                                                         
        local_tmr_voter(649)  <=    (tmr_registers(0)(649) and tmr_registers(1)(649)) or                                                             
                            (tmr_registers(1)(649) and tmr_registers(2)(649)) or                                                             
                            (tmr_registers(0)(649) and tmr_registers(2)(649));                                                               
                                                                                                                                         
        local_tmr_voter(650)  <=    (tmr_registers(0)(650) and tmr_registers(1)(650)) or                                                             
                            (tmr_registers(1)(650) and tmr_registers(2)(650)) or                                                             
                            (tmr_registers(0)(650) and tmr_registers(2)(650));                                                               
                                                                                                                                         
        local_tmr_voter(651)  <=    (tmr_registers(0)(651) and tmr_registers(1)(651)) or                                                             
                            (tmr_registers(1)(651) and tmr_registers(2)(651)) or                                                             
                            (tmr_registers(0)(651) and tmr_registers(2)(651));                                                               
                                                                                                                                         
        local_tmr_voter(652)  <=    (tmr_registers(0)(652) and tmr_registers(1)(652)) or                                                             
                            (tmr_registers(1)(652) and tmr_registers(2)(652)) or                                                             
                            (tmr_registers(0)(652) and tmr_registers(2)(652));                                                               
                                                                                                                                         
        local_tmr_voter(653)  <=    (tmr_registers(0)(653) and tmr_registers(1)(653)) or                                                             
                            (tmr_registers(1)(653) and tmr_registers(2)(653)) or                                                             
                            (tmr_registers(0)(653) and tmr_registers(2)(653));                                                               
                                                                                                                                         
        local_tmr_voter(654)  <=    (tmr_registers(0)(654) and tmr_registers(1)(654)) or                                                             
                            (tmr_registers(1)(654) and tmr_registers(2)(654)) or                                                             
                            (tmr_registers(0)(654) and tmr_registers(2)(654));                                                               
                                                                                                                                         
        local_tmr_voter(655)  <=    (tmr_registers(0)(655) and tmr_registers(1)(655)) or                                                             
                            (tmr_registers(1)(655) and tmr_registers(2)(655)) or                                                             
                            (tmr_registers(0)(655) and tmr_registers(2)(655));                                                               
                                                                                                                                         
        local_tmr_voter(656)  <=    (tmr_registers(0)(656) and tmr_registers(1)(656)) or                                                             
                            (tmr_registers(1)(656) and tmr_registers(2)(656)) or                                                             
                            (tmr_registers(0)(656) and tmr_registers(2)(656));                                                               
                                                                                                                                         
        local_tmr_voter(657)  <=    (tmr_registers(0)(657) and tmr_registers(1)(657)) or                                                             
                            (tmr_registers(1)(657) and tmr_registers(2)(657)) or                                                             
                            (tmr_registers(0)(657) and tmr_registers(2)(657));                                                               
                                                                                                                                         
        local_tmr_voter(658)  <=    (tmr_registers(0)(658) and tmr_registers(1)(658)) or                                                             
                            (tmr_registers(1)(658) and tmr_registers(2)(658)) or                                                             
                            (tmr_registers(0)(658) and tmr_registers(2)(658));                                                               
                                                                                                                                         
        local_tmr_voter(659)  <=    (tmr_registers(0)(659) and tmr_registers(1)(659)) or                                                             
                            (tmr_registers(1)(659) and tmr_registers(2)(659)) or                                                             
                            (tmr_registers(0)(659) and tmr_registers(2)(659));                                                               
                                                                                                                                         
        local_tmr_voter(660)  <=    (tmr_registers(0)(660) and tmr_registers(1)(660)) or                                                             
                            (tmr_registers(1)(660) and tmr_registers(2)(660)) or                                                             
                            (tmr_registers(0)(660) and tmr_registers(2)(660));                                                               
                                                                                                                                         
        local_tmr_voter(661)  <=    (tmr_registers(0)(661) and tmr_registers(1)(661)) or                                                             
                            (tmr_registers(1)(661) and tmr_registers(2)(661)) or                                                             
                            (tmr_registers(0)(661) and tmr_registers(2)(661));                                                               
                                                                                                                                         
        local_tmr_voter(662)  <=    (tmr_registers(0)(662) and tmr_registers(1)(662)) or                                                             
                            (tmr_registers(1)(662) and tmr_registers(2)(662)) or                                                             
                            (tmr_registers(0)(662) and tmr_registers(2)(662));                                                               
                                                                                                                                         
        local_tmr_voter(663)  <=    (tmr_registers(0)(663) and tmr_registers(1)(663)) or                                                             
                            (tmr_registers(1)(663) and tmr_registers(2)(663)) or                                                             
                            (tmr_registers(0)(663) and tmr_registers(2)(663));                                                               
                                                                                                                                         
        local_tmr_voter(664)  <=    (tmr_registers(0)(664) and tmr_registers(1)(664)) or                                                             
                            (tmr_registers(1)(664) and tmr_registers(2)(664)) or                                                             
                            (tmr_registers(0)(664) and tmr_registers(2)(664));                                                               
                                                                                                                                         
        local_tmr_voter(665)  <=    (tmr_registers(0)(665) and tmr_registers(1)(665)) or                                                             
                            (tmr_registers(1)(665) and tmr_registers(2)(665)) or                                                             
                            (tmr_registers(0)(665) and tmr_registers(2)(665));                                                               
                                                                                                                                         
        local_tmr_voter(666)  <=    (tmr_registers(0)(666) and tmr_registers(1)(666)) or                                                             
                            (tmr_registers(1)(666) and tmr_registers(2)(666)) or                                                             
                            (tmr_registers(0)(666) and tmr_registers(2)(666));                                                               
                                                                                                                                         
        local_tmr_voter(667)  <=    (tmr_registers(0)(667) and tmr_registers(1)(667)) or                                                             
                            (tmr_registers(1)(667) and tmr_registers(2)(667)) or                                                             
                            (tmr_registers(0)(667) and tmr_registers(2)(667));                                                               
                                                                                                                                         
        local_tmr_voter(668)  <=    (tmr_registers(0)(668) and tmr_registers(1)(668)) or                                                             
                            (tmr_registers(1)(668) and tmr_registers(2)(668)) or                                                             
                            (tmr_registers(0)(668) and tmr_registers(2)(668));                                                               
                                                                                                                                         
        local_tmr_voter(669)  <=    (tmr_registers(0)(669) and tmr_registers(1)(669)) or                                                             
                            (tmr_registers(1)(669) and tmr_registers(2)(669)) or                                                             
                            (tmr_registers(0)(669) and tmr_registers(2)(669));                                                               
                                                                                                                                         
        local_tmr_voter(670)  <=    (tmr_registers(0)(670) and tmr_registers(1)(670)) or                                                             
                            (tmr_registers(1)(670) and tmr_registers(2)(670)) or                                                             
                            (tmr_registers(0)(670) and tmr_registers(2)(670));                                                               
                                                                                                                                         
        local_tmr_voter(671)  <=    (tmr_registers(0)(671) and tmr_registers(1)(671)) or                                                             
                            (tmr_registers(1)(671) and tmr_registers(2)(671)) or                                                             
                            (tmr_registers(0)(671) and tmr_registers(2)(671));                                                               
                                                                                                                                         
        local_tmr_voter(672)  <=    (tmr_registers(0)(672) and tmr_registers(1)(672)) or                                                             
                            (tmr_registers(1)(672) and tmr_registers(2)(672)) or                                                             
                            (tmr_registers(0)(672) and tmr_registers(2)(672));                                                               
                                                                                                                                         
        local_tmr_voter(673)  <=    (tmr_registers(0)(673) and tmr_registers(1)(673)) or                                                             
                            (tmr_registers(1)(673) and tmr_registers(2)(673)) or                                                             
                            (tmr_registers(0)(673) and tmr_registers(2)(673));                                                               
                                                                                                                                         
        local_tmr_voter(674)  <=    (tmr_registers(0)(674) and tmr_registers(1)(674)) or                                                             
                            (tmr_registers(1)(674) and tmr_registers(2)(674)) or                                                             
                            (tmr_registers(0)(674) and tmr_registers(2)(674));                                                               
                                                                                                                                         
        local_tmr_voter(675)  <=    (tmr_registers(0)(675) and tmr_registers(1)(675)) or                                                             
                            (tmr_registers(1)(675) and tmr_registers(2)(675)) or                                                             
                            (tmr_registers(0)(675) and tmr_registers(2)(675));                                                               
                                                                                                                                         
        local_tmr_voter(676)  <=    (tmr_registers(0)(676) and tmr_registers(1)(676)) or                                                             
                            (tmr_registers(1)(676) and tmr_registers(2)(676)) or                                                             
                            (tmr_registers(0)(676) and tmr_registers(2)(676));                                                               
                                                                                                                                         
        local_tmr_voter(677)  <=    (tmr_registers(0)(677) and tmr_registers(1)(677)) or                                                             
                            (tmr_registers(1)(677) and tmr_registers(2)(677)) or                                                             
                            (tmr_registers(0)(677) and tmr_registers(2)(677));                                                               
                                                                                                                                         
        local_tmr_voter(678)  <=    (tmr_registers(0)(678) and tmr_registers(1)(678)) or                                                             
                            (tmr_registers(1)(678) and tmr_registers(2)(678)) or                                                             
                            (tmr_registers(0)(678) and tmr_registers(2)(678));                                                               
                                                                                                                                         
        local_tmr_voter(679)  <=    (tmr_registers(0)(679) and tmr_registers(1)(679)) or                                                             
                            (tmr_registers(1)(679) and tmr_registers(2)(679)) or                                                             
                            (tmr_registers(0)(679) and tmr_registers(2)(679));                                                               
                                                                                                                                         
        local_tmr_voter(680)  <=    (tmr_registers(0)(680) and tmr_registers(1)(680)) or                                                             
                            (tmr_registers(1)(680) and tmr_registers(2)(680)) or                                                             
                            (tmr_registers(0)(680) and tmr_registers(2)(680));                                                               
                                                                                                                                         
        local_tmr_voter(681)  <=    (tmr_registers(0)(681) and tmr_registers(1)(681)) or                                                             
                            (tmr_registers(1)(681) and tmr_registers(2)(681)) or                                                             
                            (tmr_registers(0)(681) and tmr_registers(2)(681));                                                               
                                                                                                                                         
        local_tmr_voter(682)  <=    (tmr_registers(0)(682) and tmr_registers(1)(682)) or                                                             
                            (tmr_registers(1)(682) and tmr_registers(2)(682)) or                                                             
                            (tmr_registers(0)(682) and tmr_registers(2)(682));                                                               
                                                                                                                                         
        local_tmr_voter(683)  <=    (tmr_registers(0)(683) and tmr_registers(1)(683)) or                                                             
                            (tmr_registers(1)(683) and tmr_registers(2)(683)) or                                                             
                            (tmr_registers(0)(683) and tmr_registers(2)(683));                                                               
                                                                                                                                         
        local_tmr_voter(684)  <=    (tmr_registers(0)(684) and tmr_registers(1)(684)) or                                                             
                            (tmr_registers(1)(684) and tmr_registers(2)(684)) or                                                             
                            (tmr_registers(0)(684) and tmr_registers(2)(684));                                                               
                                                                                                                                         
        local_tmr_voter(685)  <=    (tmr_registers(0)(685) and tmr_registers(1)(685)) or                                                             
                            (tmr_registers(1)(685) and tmr_registers(2)(685)) or                                                             
                            (tmr_registers(0)(685) and tmr_registers(2)(685));                                                               
                                                                                                                                         
        local_tmr_voter(686)  <=    (tmr_registers(0)(686) and tmr_registers(1)(686)) or                                                             
                            (tmr_registers(1)(686) and tmr_registers(2)(686)) or                                                             
                            (tmr_registers(0)(686) and tmr_registers(2)(686));                                                               
                                                                                                                                         
        local_tmr_voter(687)  <=    (tmr_registers(0)(687) and tmr_registers(1)(687)) or                                                             
                            (tmr_registers(1)(687) and tmr_registers(2)(687)) or                                                             
                            (tmr_registers(0)(687) and tmr_registers(2)(687));                                                               
                                                                                                                                         
        local_tmr_voter(688)  <=    (tmr_registers(0)(688) and tmr_registers(1)(688)) or                                                             
                            (tmr_registers(1)(688) and tmr_registers(2)(688)) or                                                             
                            (tmr_registers(0)(688) and tmr_registers(2)(688));                                                               
                                                                                                                                         
        local_tmr_voter(689)  <=    (tmr_registers(0)(689) and tmr_registers(1)(689)) or                                                             
                            (tmr_registers(1)(689) and tmr_registers(2)(689)) or                                                             
                            (tmr_registers(0)(689) and tmr_registers(2)(689));                                                               
                                                                                                                                         
        local_tmr_voter(690)  <=    (tmr_registers(0)(690) and tmr_registers(1)(690)) or                                                             
                            (tmr_registers(1)(690) and tmr_registers(2)(690)) or                                                             
                            (tmr_registers(0)(690) and tmr_registers(2)(690));                                                               
                                                                                                                                         
        local_tmr_voter(691)  <=    (tmr_registers(0)(691) and tmr_registers(1)(691)) or                                                             
                            (tmr_registers(1)(691) and tmr_registers(2)(691)) or                                                             
                            (tmr_registers(0)(691) and tmr_registers(2)(691));                                                               
                                                                                                                                         
        local_tmr_voter(692)  <=    (tmr_registers(0)(692) and tmr_registers(1)(692)) or                                                             
                            (tmr_registers(1)(692) and tmr_registers(2)(692)) or                                                             
                            (tmr_registers(0)(692) and tmr_registers(2)(692));                                                               
                                                                                                                                         
        local_tmr_voter(693)  <=    (tmr_registers(0)(693) and tmr_registers(1)(693)) or                                                             
                            (tmr_registers(1)(693) and tmr_registers(2)(693)) or                                                             
                            (tmr_registers(0)(693) and tmr_registers(2)(693));                                                               
                                                                                                                                         
        local_tmr_voter(694)  <=    (tmr_registers(0)(694) and tmr_registers(1)(694)) or                                                             
                            (tmr_registers(1)(694) and tmr_registers(2)(694)) or                                                             
                            (tmr_registers(0)(694) and tmr_registers(2)(694));                                                               
                                                                                                                                         
        local_tmr_voter(695)  <=    (tmr_registers(0)(695) and tmr_registers(1)(695)) or                                                             
                            (tmr_registers(1)(695) and tmr_registers(2)(695)) or                                                             
                            (tmr_registers(0)(695) and tmr_registers(2)(695));                                                               
                                                                                                                                         
        local_tmr_voter(696)  <=    (tmr_registers(0)(696) and tmr_registers(1)(696)) or                                                             
                            (tmr_registers(1)(696) and tmr_registers(2)(696)) or                                                             
                            (tmr_registers(0)(696) and tmr_registers(2)(696));                                                               
                                                                                                                                         
        local_tmr_voter(697)  <=    (tmr_registers(0)(697) and tmr_registers(1)(697)) or                                                             
                            (tmr_registers(1)(697) and tmr_registers(2)(697)) or                                                             
                            (tmr_registers(0)(697) and tmr_registers(2)(697));                                                               
                                                                                                                                         
        local_tmr_voter(698)  <=    (tmr_registers(0)(698) and tmr_registers(1)(698)) or                                                             
                            (tmr_registers(1)(698) and tmr_registers(2)(698)) or                                                             
                            (tmr_registers(0)(698) and tmr_registers(2)(698));                                                               
                                                                                                                                         
        local_tmr_voter(699)  <=    (tmr_registers(0)(699) and tmr_registers(1)(699)) or                                                             
                            (tmr_registers(1)(699) and tmr_registers(2)(699)) or                                                             
                            (tmr_registers(0)(699) and tmr_registers(2)(699));                                                               
                                                                                                                                         
        local_tmr_voter(700)  <=    (tmr_registers(0)(700) and tmr_registers(1)(700)) or                                                             
                            (tmr_registers(1)(700) and tmr_registers(2)(700)) or                                                             
                            (tmr_registers(0)(700) and tmr_registers(2)(700));                                                               
                                                                                                                                         
        local_tmr_voter(701)  <=    (tmr_registers(0)(701) and tmr_registers(1)(701)) or                                                             
                            (tmr_registers(1)(701) and tmr_registers(2)(701)) or                                                             
                            (tmr_registers(0)(701) and tmr_registers(2)(701));                                                               
                                                                                                                                         
        local_tmr_voter(702)  <=    (tmr_registers(0)(702) and tmr_registers(1)(702)) or                                                             
                            (tmr_registers(1)(702) and tmr_registers(2)(702)) or                                                             
                            (tmr_registers(0)(702) and tmr_registers(2)(702));                                                               
                                                                                                                                         
        local_tmr_voter(703)  <=    (tmr_registers(0)(703) and tmr_registers(1)(703)) or                                                             
                            (tmr_registers(1)(703) and tmr_registers(2)(703)) or                                                             
                            (tmr_registers(0)(703) and tmr_registers(2)(703));                                                               
                                                                                                                                         
        local_tmr_voter(704)  <=    (tmr_registers(0)(704) and tmr_registers(1)(704)) or                                                             
                            (tmr_registers(1)(704) and tmr_registers(2)(704)) or                                                             
                            (tmr_registers(0)(704) and tmr_registers(2)(704));                                                               
                                                                                                                                         
        local_tmr_voter(705)  <=    (tmr_registers(0)(705) and tmr_registers(1)(705)) or                                                             
                            (tmr_registers(1)(705) and tmr_registers(2)(705)) or                                                             
                            (tmr_registers(0)(705) and tmr_registers(2)(705));                                                               
                                                                                                                                         
        local_tmr_voter(706)  <=    (tmr_registers(0)(706) and tmr_registers(1)(706)) or                                                             
                            (tmr_registers(1)(706) and tmr_registers(2)(706)) or                                                             
                            (tmr_registers(0)(706) and tmr_registers(2)(706));                                                               
                                                                                                                                         
        local_tmr_voter(707)  <=    (tmr_registers(0)(707) and tmr_registers(1)(707)) or                                                             
                            (tmr_registers(1)(707) and tmr_registers(2)(707)) or                                                             
                            (tmr_registers(0)(707) and tmr_registers(2)(707));                                                               
                                                                                                                                         
        local_tmr_voter(708)  <=    (tmr_registers(0)(708) and tmr_registers(1)(708)) or                                                             
                            (tmr_registers(1)(708) and tmr_registers(2)(708)) or                                                             
                            (tmr_registers(0)(708) and tmr_registers(2)(708));                                                               
                                                                                                                                         
        local_tmr_voter(709)  <=    (tmr_registers(0)(709) and tmr_registers(1)(709)) or                                                             
                            (tmr_registers(1)(709) and tmr_registers(2)(709)) or                                                             
                            (tmr_registers(0)(709) and tmr_registers(2)(709));                                                               
                                                                                                                                         
        local_tmr_voter(710)  <=    (tmr_registers(0)(710) and tmr_registers(1)(710)) or                                                             
                            (tmr_registers(1)(710) and tmr_registers(2)(710)) or                                                             
                            (tmr_registers(0)(710) and tmr_registers(2)(710));                                                               
                                                                                                                                         
        local_tmr_voter(711)  <=    (tmr_registers(0)(711) and tmr_registers(1)(711)) or                                                             
                            (tmr_registers(1)(711) and tmr_registers(2)(711)) or                                                             
                            (tmr_registers(0)(711) and tmr_registers(2)(711));                                                               
                                                                                                                                         
        local_tmr_voter(712)  <=    (tmr_registers(0)(712) and tmr_registers(1)(712)) or                                                             
                            (tmr_registers(1)(712) and tmr_registers(2)(712)) or                                                             
                            (tmr_registers(0)(712) and tmr_registers(2)(712));                                                               
                                                                                                                                         
        local_tmr_voter(713)  <=    (tmr_registers(0)(713) and tmr_registers(1)(713)) or                                                             
                            (tmr_registers(1)(713) and tmr_registers(2)(713)) or                                                             
                            (tmr_registers(0)(713) and tmr_registers(2)(713));                                                               
                                                                                                                                         
        local_tmr_voter(714)  <=    (tmr_registers(0)(714) and tmr_registers(1)(714)) or                                                             
                            (tmr_registers(1)(714) and tmr_registers(2)(714)) or                                                             
                            (tmr_registers(0)(714) and tmr_registers(2)(714));                                                               
                                                                                                                                         
        local_tmr_voter(715)  <=    (tmr_registers(0)(715) and tmr_registers(1)(715)) or                                                             
                            (tmr_registers(1)(715) and tmr_registers(2)(715)) or                                                             
                            (tmr_registers(0)(715) and tmr_registers(2)(715));                                                               
                                                                                                                                         
        local_tmr_voter(716)  <=    (tmr_registers(0)(716) and tmr_registers(1)(716)) or                                                             
                            (tmr_registers(1)(716) and tmr_registers(2)(716)) or                                                             
                            (tmr_registers(0)(716) and tmr_registers(2)(716));                                                               
                                                                                                                                         
        local_tmr_voter(717)  <=    (tmr_registers(0)(717) and tmr_registers(1)(717)) or                                                             
                            (tmr_registers(1)(717) and tmr_registers(2)(717)) or                                                             
                            (tmr_registers(0)(717) and tmr_registers(2)(717));                                                               
                                                                                                                                         
        local_tmr_voter(718)  <=    (tmr_registers(0)(718) and tmr_registers(1)(718)) or                                                             
                            (tmr_registers(1)(718) and tmr_registers(2)(718)) or                                                             
                            (tmr_registers(0)(718) and tmr_registers(2)(718));                                                               
                                                                                                                                         
        local_tmr_voter(719)  <=    (tmr_registers(0)(719) and tmr_registers(1)(719)) or                                                             
                            (tmr_registers(1)(719) and tmr_registers(2)(719)) or                                                             
                            (tmr_registers(0)(719) and tmr_registers(2)(719));                                                               
                                                                                                                                         
        local_tmr_voter(720)  <=    (tmr_registers(0)(720) and tmr_registers(1)(720)) or                                                             
                            (tmr_registers(1)(720) and tmr_registers(2)(720)) or                                                             
                            (tmr_registers(0)(720) and tmr_registers(2)(720));                                                               
                                                                                                                                         
        local_tmr_voter(721)  <=    (tmr_registers(0)(721) and tmr_registers(1)(721)) or                                                             
                            (tmr_registers(1)(721) and tmr_registers(2)(721)) or                                                             
                            (tmr_registers(0)(721) and tmr_registers(2)(721));                                                               
                                                                                                                                         
        local_tmr_voter(722)  <=    (tmr_registers(0)(722) and tmr_registers(1)(722)) or                                                             
                            (tmr_registers(1)(722) and tmr_registers(2)(722)) or                                                             
                            (tmr_registers(0)(722) and tmr_registers(2)(722));                                                               
                                                                                                                                         
        local_tmr_voter(723)  <=    (tmr_registers(0)(723) and tmr_registers(1)(723)) or                                                             
                            (tmr_registers(1)(723) and tmr_registers(2)(723)) or                                                             
                            (tmr_registers(0)(723) and tmr_registers(2)(723));                                                               
                                                                                                                                         
        local_tmr_voter(724)  <=    (tmr_registers(0)(724) and tmr_registers(1)(724)) or                                                             
                            (tmr_registers(1)(724) and tmr_registers(2)(724)) or                                                             
                            (tmr_registers(0)(724) and tmr_registers(2)(724));                                                               
                                                                                                                                         
        local_tmr_voter(725)  <=    (tmr_registers(0)(725) and tmr_registers(1)(725)) or                                                             
                            (tmr_registers(1)(725) and tmr_registers(2)(725)) or                                                             
                            (tmr_registers(0)(725) and tmr_registers(2)(725));                                                               
                                                                                                                                         
        local_tmr_voter(726)  <=    (tmr_registers(0)(726) and tmr_registers(1)(726)) or                                                             
                            (tmr_registers(1)(726) and tmr_registers(2)(726)) or                                                             
                            (tmr_registers(0)(726) and tmr_registers(2)(726));                                                               
                                                                                                                                         
        local_tmr_voter(727)  <=    (tmr_registers(0)(727) and tmr_registers(1)(727)) or                                                             
                            (tmr_registers(1)(727) and tmr_registers(2)(727)) or                                                             
                            (tmr_registers(0)(727) and tmr_registers(2)(727));                                                               
                                                                                                                                         
        local_tmr_voter(728)  <=    (tmr_registers(0)(728) and tmr_registers(1)(728)) or                                                             
                            (tmr_registers(1)(728) and tmr_registers(2)(728)) or                                                             
                            (tmr_registers(0)(728) and tmr_registers(2)(728));                                                               
                                                                                                                                         
        local_tmr_voter(729)  <=    (tmr_registers(0)(729) and tmr_registers(1)(729)) or                                                             
                            (tmr_registers(1)(729) and tmr_registers(2)(729)) or                                                             
                            (tmr_registers(0)(729) and tmr_registers(2)(729));                                                               
                                                                                                                                         
        local_tmr_voter(730)  <=    (tmr_registers(0)(730) and tmr_registers(1)(730)) or                                                             
                            (tmr_registers(1)(730) and tmr_registers(2)(730)) or                                                             
                            (tmr_registers(0)(730) and tmr_registers(2)(730));                                                               
                                                                                                                                         
        local_tmr_voter(731)  <=    (tmr_registers(0)(731) and tmr_registers(1)(731)) or                                                             
                            (tmr_registers(1)(731) and tmr_registers(2)(731)) or                                                             
                            (tmr_registers(0)(731) and tmr_registers(2)(731));                                                               
                                                                                                                                         
        local_tmr_voter(732)  <=    (tmr_registers(0)(732) and tmr_registers(1)(732)) or                                                             
                            (tmr_registers(1)(732) and tmr_registers(2)(732)) or                                                             
                            (tmr_registers(0)(732) and tmr_registers(2)(732));                                                               
                                                                                                                                         
        local_tmr_voter(733)  <=    (tmr_registers(0)(733) and tmr_registers(1)(733)) or                                                             
                            (tmr_registers(1)(733) and tmr_registers(2)(733)) or                                                             
                            (tmr_registers(0)(733) and tmr_registers(2)(733));                                                               
                                                                                                                                         
        local_tmr_voter(734)  <=    (tmr_registers(0)(734) and tmr_registers(1)(734)) or                                                             
                            (tmr_registers(1)(734) and tmr_registers(2)(734)) or                                                             
                            (tmr_registers(0)(734) and tmr_registers(2)(734));                                                               
                                                                                                                                         
        local_tmr_voter(735)  <=    (tmr_registers(0)(735) and tmr_registers(1)(735)) or                                                             
                            (tmr_registers(1)(735) and tmr_registers(2)(735)) or                                                             
                            (tmr_registers(0)(735) and tmr_registers(2)(735));                                                               
                                                                                                                                         
        local_tmr_voter(736)  <=    (tmr_registers(0)(736) and tmr_registers(1)(736)) or                                                             
                            (tmr_registers(1)(736) and tmr_registers(2)(736)) or                                                             
                            (tmr_registers(0)(736) and tmr_registers(2)(736));                                                               
                                                                                                                                         
        local_tmr_voter(737)  <=    (tmr_registers(0)(737) and tmr_registers(1)(737)) or                                                             
                            (tmr_registers(1)(737) and tmr_registers(2)(737)) or                                                             
                            (tmr_registers(0)(737) and tmr_registers(2)(737));                                                               
                                                                                                                                         
        local_tmr_voter(738)  <=    (tmr_registers(0)(738) and tmr_registers(1)(738)) or                                                             
                            (tmr_registers(1)(738) and tmr_registers(2)(738)) or                                                             
                            (tmr_registers(0)(738) and tmr_registers(2)(738));                                                               
                                                                                                                                         
        local_tmr_voter(739)  <=    (tmr_registers(0)(739) and tmr_registers(1)(739)) or                                                             
                            (tmr_registers(1)(739) and tmr_registers(2)(739)) or                                                             
                            (tmr_registers(0)(739) and tmr_registers(2)(739));                                                               
                                                                                                                                         
        local_tmr_voter(740)  <=    (tmr_registers(0)(740) and tmr_registers(1)(740)) or                                                             
                            (tmr_registers(1)(740) and tmr_registers(2)(740)) or                                                             
                            (tmr_registers(0)(740) and tmr_registers(2)(740));                                                               
                                                                                                                                         
        local_tmr_voter(741)  <=    (tmr_registers(0)(741) and tmr_registers(1)(741)) or                                                             
                            (tmr_registers(1)(741) and tmr_registers(2)(741)) or                                                             
                            (tmr_registers(0)(741) and tmr_registers(2)(741));                                                               
                                                                                                                                         
        local_tmr_voter(742)  <=    (tmr_registers(0)(742) and tmr_registers(1)(742)) or                                                             
                            (tmr_registers(1)(742) and tmr_registers(2)(742)) or                                                             
                            (tmr_registers(0)(742) and tmr_registers(2)(742));                                                               
                                                                                                                                         
        local_tmr_voter(743)  <=    (tmr_registers(0)(743) and tmr_registers(1)(743)) or                                                             
                            (tmr_registers(1)(743) and tmr_registers(2)(743)) or                                                             
                            (tmr_registers(0)(743) and tmr_registers(2)(743));                                                               
                                                                                                                                         
        local_tmr_voter(744)  <=    (tmr_registers(0)(744) and tmr_registers(1)(744)) or                                                             
                            (tmr_registers(1)(744) and tmr_registers(2)(744)) or                                                             
                            (tmr_registers(0)(744) and tmr_registers(2)(744));                                                               
                                                                                                                                         
        local_tmr_voter(745)  <=    (tmr_registers(0)(745) and tmr_registers(1)(745)) or                                                             
                            (tmr_registers(1)(745) and tmr_registers(2)(745)) or                                                             
                            (tmr_registers(0)(745) and tmr_registers(2)(745));                                                               
                                                                                                                                         
        local_tmr_voter(746)  <=    (tmr_registers(0)(746) and tmr_registers(1)(746)) or                                                             
                            (tmr_registers(1)(746) and tmr_registers(2)(746)) or                                                             
                            (tmr_registers(0)(746) and tmr_registers(2)(746));                                                               
                                                                                                                                         
        local_tmr_voter(747)  <=    (tmr_registers(0)(747) and tmr_registers(1)(747)) or                                                             
                            (tmr_registers(1)(747) and tmr_registers(2)(747)) or                                                             
                            (tmr_registers(0)(747) and tmr_registers(2)(747));                                                               
                                                                                                                                         
        local_tmr_voter(748)  <=    (tmr_registers(0)(748) and tmr_registers(1)(748)) or                                                             
                            (tmr_registers(1)(748) and tmr_registers(2)(748)) or                                                             
                            (tmr_registers(0)(748) and tmr_registers(2)(748));                                                               
                                                                                                                                         
        local_tmr_voter(749)  <=    (tmr_registers(0)(749) and tmr_registers(1)(749)) or                                                             
                            (tmr_registers(1)(749) and tmr_registers(2)(749)) or                                                             
                            (tmr_registers(0)(749) and tmr_registers(2)(749));                                                               
                                                                                                                                         
        local_tmr_voter(750)  <=    (tmr_registers(0)(750) and tmr_registers(1)(750)) or                                                             
                            (tmr_registers(1)(750) and tmr_registers(2)(750)) or                                                             
                            (tmr_registers(0)(750) and tmr_registers(2)(750));                                                               
                                                                                                                                         
        local_tmr_voter(751)  <=    (tmr_registers(0)(751) and tmr_registers(1)(751)) or                                                             
                            (tmr_registers(1)(751) and tmr_registers(2)(751)) or                                                             
                            (tmr_registers(0)(751) and tmr_registers(2)(751));                                                               
                                                                                                                                         
        local_tmr_voter(752)  <=    (tmr_registers(0)(752) and tmr_registers(1)(752)) or                                                             
                            (tmr_registers(1)(752) and tmr_registers(2)(752)) or                                                             
                            (tmr_registers(0)(752) and tmr_registers(2)(752));                                                               
                                                                                                                                         
        local_tmr_voter(753)  <=    (tmr_registers(0)(753) and tmr_registers(1)(753)) or                                                             
                            (tmr_registers(1)(753) and tmr_registers(2)(753)) or                                                             
                            (tmr_registers(0)(753) and tmr_registers(2)(753));                                                               
                                                                                                                                         
        local_tmr_voter(754)  <=    (tmr_registers(0)(754) and tmr_registers(1)(754)) or                                                             
                            (tmr_registers(1)(754) and tmr_registers(2)(754)) or                                                             
                            (tmr_registers(0)(754) and tmr_registers(2)(754));                                                               
                                                                                                                                         
        local_tmr_voter(755)  <=    (tmr_registers(0)(755) and tmr_registers(1)(755)) or                                                             
                            (tmr_registers(1)(755) and tmr_registers(2)(755)) or                                                             
                            (tmr_registers(0)(755) and tmr_registers(2)(755));                                                               
                                                                                                                                         
        local_tmr_voter(756)  <=    (tmr_registers(0)(756) and tmr_registers(1)(756)) or                                                             
                            (tmr_registers(1)(756) and tmr_registers(2)(756)) or                                                             
                            (tmr_registers(0)(756) and tmr_registers(2)(756));                                                               
                                                                                                                                         
        local_tmr_voter(757)  <=    (tmr_registers(0)(757) and tmr_registers(1)(757)) or                                                             
                            (tmr_registers(1)(757) and tmr_registers(2)(757)) or                                                             
                            (tmr_registers(0)(757) and tmr_registers(2)(757));                                                               
                                                                                                                                         
        local_tmr_voter(758)  <=    (tmr_registers(0)(758) and tmr_registers(1)(758)) or                                                             
                            (tmr_registers(1)(758) and tmr_registers(2)(758)) or                                                             
                            (tmr_registers(0)(758) and tmr_registers(2)(758));                                                               
                                                                                                                                         
        local_tmr_voter(759)  <=    (tmr_registers(0)(759) and tmr_registers(1)(759)) or                                                             
                            (tmr_registers(1)(759) and tmr_registers(2)(759)) or                                                             
                            (tmr_registers(0)(759) and tmr_registers(2)(759));                                                               
                                                                                                                                         
        local_tmr_voter(760)  <=    (tmr_registers(0)(760) and tmr_registers(1)(760)) or                                                             
                            (tmr_registers(1)(760) and tmr_registers(2)(760)) or                                                             
                            (tmr_registers(0)(760) and tmr_registers(2)(760));                                                               
                                                                                                                                         
        local_tmr_voter(761)  <=    (tmr_registers(0)(761) and tmr_registers(1)(761)) or                                                             
                            (tmr_registers(1)(761) and tmr_registers(2)(761)) or                                                             
                            (tmr_registers(0)(761) and tmr_registers(2)(761));                                                               
                                                                                                                                         
        local_tmr_voter(762)  <=    (tmr_registers(0)(762) and tmr_registers(1)(762)) or                                                             
                            (tmr_registers(1)(762) and tmr_registers(2)(762)) or                                                             
                            (tmr_registers(0)(762) and tmr_registers(2)(762));                                                               
                                                                                                                                         
        local_tmr_voter(763)  <=    (tmr_registers(0)(763) and tmr_registers(1)(763)) or                                                             
                            (tmr_registers(1)(763) and tmr_registers(2)(763)) or                                                             
                            (tmr_registers(0)(763) and tmr_registers(2)(763));                                                               
                                                                                                                                         
        local_tmr_voter(764)  <=    (tmr_registers(0)(764) and tmr_registers(1)(764)) or                                                             
                            (tmr_registers(1)(764) and tmr_registers(2)(764)) or                                                             
                            (tmr_registers(0)(764) and tmr_registers(2)(764));                                                               
                                                                                                                                         
        local_tmr_voter(765)  <=    (tmr_registers(0)(765) and tmr_registers(1)(765)) or                                                             
                            (tmr_registers(1)(765) and tmr_registers(2)(765)) or                                                             
                            (tmr_registers(0)(765) and tmr_registers(2)(765));                                                               
                                                                                                                                         
        local_tmr_voter(766)  <=    (tmr_registers(0)(766) and tmr_registers(1)(766)) or                                                             
                            (tmr_registers(1)(766) and tmr_registers(2)(766)) or                                                             
                            (tmr_registers(0)(766) and tmr_registers(2)(766));                                                               
                                                                                                                                         
        local_tmr_voter(767)  <=    (tmr_registers(0)(767) and tmr_registers(1)(767)) or                                                             
                            (tmr_registers(1)(767) and tmr_registers(2)(767)) or                                                             
                            (tmr_registers(0)(767) and tmr_registers(2)(767));                                                               
                                                                                                                                         
        local_tmr_voter(768)  <=    (tmr_registers(0)(768) and tmr_registers(1)(768)) or                                                             
                            (tmr_registers(1)(768) and tmr_registers(2)(768)) or                                                             
                            (tmr_registers(0)(768) and tmr_registers(2)(768));                                                               
                                                                                                                                         
        local_tmr_voter(769)  <=    (tmr_registers(0)(769) and tmr_registers(1)(769)) or                                                             
                            (tmr_registers(1)(769) and tmr_registers(2)(769)) or                                                             
                            (tmr_registers(0)(769) and tmr_registers(2)(769));                                                               
                                                                                                                                         
        local_tmr_voter(770)  <=    (tmr_registers(0)(770) and tmr_registers(1)(770)) or                                                             
                            (tmr_registers(1)(770) and tmr_registers(2)(770)) or                                                             
                            (tmr_registers(0)(770) and tmr_registers(2)(770));                                                               
                                                                                                                                         
        local_tmr_voter(771)  <=    (tmr_registers(0)(771) and tmr_registers(1)(771)) or                                                             
                            (tmr_registers(1)(771) and tmr_registers(2)(771)) or                                                             
                            (tmr_registers(0)(771) and tmr_registers(2)(771));                                                               
                                                                                                                                         
        local_tmr_voter(772)  <=    (tmr_registers(0)(772) and tmr_registers(1)(772)) or                                                             
                            (tmr_registers(1)(772) and tmr_registers(2)(772)) or                                                             
                            (tmr_registers(0)(772) and tmr_registers(2)(772));                                                               
                                                                                                                                         
        local_tmr_voter(773)  <=    (tmr_registers(0)(773) and tmr_registers(1)(773)) or                                                             
                            (tmr_registers(1)(773) and tmr_registers(2)(773)) or                                                             
                            (tmr_registers(0)(773) and tmr_registers(2)(773));                                                               
                                                                                                                                         
        local_tmr_voter(774)  <=    (tmr_registers(0)(774) and tmr_registers(1)(774)) or                                                             
                            (tmr_registers(1)(774) and tmr_registers(2)(774)) or                                                             
                            (tmr_registers(0)(774) and tmr_registers(2)(774));                                                               
                                                                                                                                         
        local_tmr_voter(775)  <=    (tmr_registers(0)(775) and tmr_registers(1)(775)) or                                                             
                            (tmr_registers(1)(775) and tmr_registers(2)(775)) or                                                             
                            (tmr_registers(0)(775) and tmr_registers(2)(775));                                                               
                                                                                                                                         
        local_tmr_voter(776)  <=    (tmr_registers(0)(776) and tmr_registers(1)(776)) or                                                             
                            (tmr_registers(1)(776) and tmr_registers(2)(776)) or                                                             
                            (tmr_registers(0)(776) and tmr_registers(2)(776));                                                               
                                                                                                                                         
        local_tmr_voter(777)  <=    (tmr_registers(0)(777) and tmr_registers(1)(777)) or                                                             
                            (tmr_registers(1)(777) and tmr_registers(2)(777)) or                                                             
                            (tmr_registers(0)(777) and tmr_registers(2)(777));                                                               
                                                                                                                                         
        local_tmr_voter(778)  <=    (tmr_registers(0)(778) and tmr_registers(1)(778)) or                                                             
                            (tmr_registers(1)(778) and tmr_registers(2)(778)) or                                                             
                            (tmr_registers(0)(778) and tmr_registers(2)(778));                                                               
                                                                                                                                         
        local_tmr_voter(779)  <=    (tmr_registers(0)(779) and tmr_registers(1)(779)) or                                                             
                            (tmr_registers(1)(779) and tmr_registers(2)(779)) or                                                             
                            (tmr_registers(0)(779) and tmr_registers(2)(779));                                                               
                                                                                                                                         
        local_tmr_voter(780)  <=    (tmr_registers(0)(780) and tmr_registers(1)(780)) or                                                             
                            (tmr_registers(1)(780) and tmr_registers(2)(780)) or                                                             
                            (tmr_registers(0)(780) and tmr_registers(2)(780));                                                               
                                                                                                                                         
        local_tmr_voter(781)  <=    (tmr_registers(0)(781) and tmr_registers(1)(781)) or                                                             
                            (tmr_registers(1)(781) and tmr_registers(2)(781)) or                                                             
                            (tmr_registers(0)(781) and tmr_registers(2)(781));                                                               
                                                                                                                                         
        local_tmr_voter(782)  <=    (tmr_registers(0)(782) and tmr_registers(1)(782)) or                                                             
                            (tmr_registers(1)(782) and tmr_registers(2)(782)) or                                                             
                            (tmr_registers(0)(782) and tmr_registers(2)(782));                                                               
                                                                                                                                         
        local_tmr_voter(783)  <=    (tmr_registers(0)(783) and tmr_registers(1)(783)) or                                                             
                            (tmr_registers(1)(783) and tmr_registers(2)(783)) or                                                             
                            (tmr_registers(0)(783) and tmr_registers(2)(783));                                                               
                                                                                                                                         
        local_tmr_voter(784)  <=    (tmr_registers(0)(784) and tmr_registers(1)(784)) or                                                             
                            (tmr_registers(1)(784) and tmr_registers(2)(784)) or                                                             
                            (tmr_registers(0)(784) and tmr_registers(2)(784));                                                               
                                                                                                                                         
        local_tmr_voter(785)  <=    (tmr_registers(0)(785) and tmr_registers(1)(785)) or                                                             
                            (tmr_registers(1)(785) and tmr_registers(2)(785)) or                                                             
                            (tmr_registers(0)(785) and tmr_registers(2)(785));                                                               
                                                                                                                                         
        local_tmr_voter(786)  <=    (tmr_registers(0)(786) and tmr_registers(1)(786)) or                                                             
                            (tmr_registers(1)(786) and tmr_registers(2)(786)) or                                                             
                            (tmr_registers(0)(786) and tmr_registers(2)(786));                                                               
                                                                                                                                         
        local_tmr_voter(787)  <=    (tmr_registers(0)(787) and tmr_registers(1)(787)) or                                                             
                            (tmr_registers(1)(787) and tmr_registers(2)(787)) or                                                             
                            (tmr_registers(0)(787) and tmr_registers(2)(787));                                                               
                                                                                                                                         
        local_tmr_voter(788)  <=    (tmr_registers(0)(788) and tmr_registers(1)(788)) or                                                             
                            (tmr_registers(1)(788) and tmr_registers(2)(788)) or                                                             
                            (tmr_registers(0)(788) and tmr_registers(2)(788));                                                               
                                                                                                                                         
        local_tmr_voter(789)  <=    (tmr_registers(0)(789) and tmr_registers(1)(789)) or                                                             
                            (tmr_registers(1)(789) and tmr_registers(2)(789)) or                                                             
                            (tmr_registers(0)(789) and tmr_registers(2)(789));                                                               
                                                                                                                                         
        local_tmr_voter(790)  <=    (tmr_registers(0)(790) and tmr_registers(1)(790)) or                                                             
                            (tmr_registers(1)(790) and tmr_registers(2)(790)) or                                                             
                            (tmr_registers(0)(790) and tmr_registers(2)(790));                                                               
                                                                                                                                         
        local_tmr_voter(791)  <=    (tmr_registers(0)(791) and tmr_registers(1)(791)) or                                                             
                            (tmr_registers(1)(791) and tmr_registers(2)(791)) or                                                             
                            (tmr_registers(0)(791) and tmr_registers(2)(791));                                                               
                                                                                                                                         
        local_tmr_voter(792)  <=    (tmr_registers(0)(792) and tmr_registers(1)(792)) or                                                             
                            (tmr_registers(1)(792) and tmr_registers(2)(792)) or                                                             
                            (tmr_registers(0)(792) and tmr_registers(2)(792));                                                               
                                                                                                                                         
        local_tmr_voter(793)  <=    (tmr_registers(0)(793) and tmr_registers(1)(793)) or                                                             
                            (tmr_registers(1)(793) and tmr_registers(2)(793)) or                                                             
                            (tmr_registers(0)(793) and tmr_registers(2)(793));                                                               
                                                                                                                                         
        local_tmr_voter(794)  <=    (tmr_registers(0)(794) and tmr_registers(1)(794)) or                                                             
                            (tmr_registers(1)(794) and tmr_registers(2)(794)) or                                                             
                            (tmr_registers(0)(794) and tmr_registers(2)(794));                                                               
                                                                                                                                         
        local_tmr_voter(795)  <=    (tmr_registers(0)(795) and tmr_registers(1)(795)) or                                                             
                            (tmr_registers(1)(795) and tmr_registers(2)(795)) or                                                             
                            (tmr_registers(0)(795) and tmr_registers(2)(795));                                                               
                                                                                                                                         
        local_tmr_voter(796)  <=    (tmr_registers(0)(796) and tmr_registers(1)(796)) or                                                             
                            (tmr_registers(1)(796) and tmr_registers(2)(796)) or                                                             
                            (tmr_registers(0)(796) and tmr_registers(2)(796));                                                               
                                                                                                                                         
        local_tmr_voter(797)  <=    (tmr_registers(0)(797) and tmr_registers(1)(797)) or                                                             
                            (tmr_registers(1)(797) and tmr_registers(2)(797)) or                                                             
                            (tmr_registers(0)(797) and tmr_registers(2)(797));                                                               
                                                                                                                                         
        local_tmr_voter(798)  <=    (tmr_registers(0)(798) and tmr_registers(1)(798)) or                                                             
                            (tmr_registers(1)(798) and tmr_registers(2)(798)) or                                                             
                            (tmr_registers(0)(798) and tmr_registers(2)(798));                                                               
                                                                                                                                         
        local_tmr_voter(799)  <=    (tmr_registers(0)(799) and tmr_registers(1)(799)) or                                                             
                            (tmr_registers(1)(799) and tmr_registers(2)(799)) or                                                             
                            (tmr_registers(0)(799) and tmr_registers(2)(799));                                                               
                                                                                                                                         
        local_tmr_voter(800)  <=    (tmr_registers(0)(800) and tmr_registers(1)(800)) or                                                             
                            (tmr_registers(1)(800) and tmr_registers(2)(800)) or                                                             
                            (tmr_registers(0)(800) and tmr_registers(2)(800));                                                               
                                                                                                                                         
        local_tmr_voter(801)  <=    (tmr_registers(0)(801) and tmr_registers(1)(801)) or                                                             
                            (tmr_registers(1)(801) and tmr_registers(2)(801)) or                                                             
                            (tmr_registers(0)(801) and tmr_registers(2)(801));                                                               
                                                                                                                                         
        local_tmr_voter(802)  <=    (tmr_registers(0)(802) and tmr_registers(1)(802)) or                                                             
                            (tmr_registers(1)(802) and tmr_registers(2)(802)) or                                                             
                            (tmr_registers(0)(802) and tmr_registers(2)(802));                                                               
                                                                                                                                         
        local_tmr_voter(803)  <=    (tmr_registers(0)(803) and tmr_registers(1)(803)) or                                                             
                            (tmr_registers(1)(803) and tmr_registers(2)(803)) or                                                             
                            (tmr_registers(0)(803) and tmr_registers(2)(803));                                                               
                                                                                                                                         
        local_tmr_voter(804)  <=    (tmr_registers(0)(804) and tmr_registers(1)(804)) or                                                             
                            (tmr_registers(1)(804) and tmr_registers(2)(804)) or                                                             
                            (tmr_registers(0)(804) and tmr_registers(2)(804));                                                               
                                                                                                                                         
        local_tmr_voter(805)  <=    (tmr_registers(0)(805) and tmr_registers(1)(805)) or                                                             
                            (tmr_registers(1)(805) and tmr_registers(2)(805)) or                                                             
                            (tmr_registers(0)(805) and tmr_registers(2)(805));                                                               
                                                                                                                                         
        local_tmr_voter(806)  <=    (tmr_registers(0)(806) and tmr_registers(1)(806)) or                                                             
                            (tmr_registers(1)(806) and tmr_registers(2)(806)) or                                                             
                            (tmr_registers(0)(806) and tmr_registers(2)(806));                                                               
                                                                                                                                         
        local_tmr_voter(807)  <=    (tmr_registers(0)(807) and tmr_registers(1)(807)) or                                                             
                            (tmr_registers(1)(807) and tmr_registers(2)(807)) or                                                             
                            (tmr_registers(0)(807) and tmr_registers(2)(807));                                                               
                                                                                                                                         
        local_tmr_voter(808)  <=    (tmr_registers(0)(808) and tmr_registers(1)(808)) or                                                             
                            (tmr_registers(1)(808) and tmr_registers(2)(808)) or                                                             
                            (tmr_registers(0)(808) and tmr_registers(2)(808));                                                               
                                                                                                                                         
        local_tmr_voter(809)  <=    (tmr_registers(0)(809) and tmr_registers(1)(809)) or                                                             
                            (tmr_registers(1)(809) and tmr_registers(2)(809)) or                                                             
                            (tmr_registers(0)(809) and tmr_registers(2)(809));                                                               
                                                                                                                                         
        local_tmr_voter(810)  <=    (tmr_registers(0)(810) and tmr_registers(1)(810)) or                                                             
                            (tmr_registers(1)(810) and tmr_registers(2)(810)) or                                                             
                            (tmr_registers(0)(810) and tmr_registers(2)(810));                                                               
                                                                                                                                         
        local_tmr_voter(811)  <=    (tmr_registers(0)(811) and tmr_registers(1)(811)) or                                                             
                            (tmr_registers(1)(811) and tmr_registers(2)(811)) or                                                             
                            (tmr_registers(0)(811) and tmr_registers(2)(811));                                                               
                                                                                                                                         
        local_tmr_voter(812)  <=    (tmr_registers(0)(812) and tmr_registers(1)(812)) or                                                             
                            (tmr_registers(1)(812) and tmr_registers(2)(812)) or                                                             
                            (tmr_registers(0)(812) and tmr_registers(2)(812));                                                               
                                                                                                                                         
        local_tmr_voter(813)  <=    (tmr_registers(0)(813) and tmr_registers(1)(813)) or                                                             
                            (tmr_registers(1)(813) and tmr_registers(2)(813)) or                                                             
                            (tmr_registers(0)(813) and tmr_registers(2)(813));                                                               
                                                                                                                                         
        local_tmr_voter(814)  <=    (tmr_registers(0)(814) and tmr_registers(1)(814)) or                                                             
                            (tmr_registers(1)(814) and tmr_registers(2)(814)) or                                                             
                            (tmr_registers(0)(814) and tmr_registers(2)(814));                                                               
                                                                                                                                         
        local_tmr_voter(815)  <=    (tmr_registers(0)(815) and tmr_registers(1)(815)) or                                                             
                            (tmr_registers(1)(815) and tmr_registers(2)(815)) or                                                             
                            (tmr_registers(0)(815) and tmr_registers(2)(815));                                                               
                                                                                                                                         
        local_tmr_voter(816)  <=    (tmr_registers(0)(816) and tmr_registers(1)(816)) or                                                             
                            (tmr_registers(1)(816) and tmr_registers(2)(816)) or                                                             
                            (tmr_registers(0)(816) and tmr_registers(2)(816));                                                               
                                                                                                                                         
        local_tmr_voter(817)  <=    (tmr_registers(0)(817) and tmr_registers(1)(817)) or                                                             
                            (tmr_registers(1)(817) and tmr_registers(2)(817)) or                                                             
                            (tmr_registers(0)(817) and tmr_registers(2)(817));                                                               
                                                                                                                                         
        local_tmr_voter(818)  <=    (tmr_registers(0)(818) and tmr_registers(1)(818)) or                                                             
                            (tmr_registers(1)(818) and tmr_registers(2)(818)) or                                                             
                            (tmr_registers(0)(818) and tmr_registers(2)(818));                                                               
                                                                                                                                         
        local_tmr_voter(819)  <=    (tmr_registers(0)(819) and tmr_registers(1)(819)) or                                                             
                            (tmr_registers(1)(819) and tmr_registers(2)(819)) or                                                             
                            (tmr_registers(0)(819) and tmr_registers(2)(819));                                                               
                                                                                                                                         
        local_tmr_voter(820)  <=    (tmr_registers(0)(820) and tmr_registers(1)(820)) or                                                             
                            (tmr_registers(1)(820) and tmr_registers(2)(820)) or                                                             
                            (tmr_registers(0)(820) and tmr_registers(2)(820));                                                               
                                                                                                                                         
        local_tmr_voter(821)  <=    (tmr_registers(0)(821) and tmr_registers(1)(821)) or                                                             
                            (tmr_registers(1)(821) and tmr_registers(2)(821)) or                                                             
                            (tmr_registers(0)(821) and tmr_registers(2)(821));                                                               
                                                                                                                                         
        local_tmr_voter(822)  <=    (tmr_registers(0)(822) and tmr_registers(1)(822)) or                                                             
                            (tmr_registers(1)(822) and tmr_registers(2)(822)) or                                                             
                            (tmr_registers(0)(822) and tmr_registers(2)(822));                                                               
                                                                                                                                         
        local_tmr_voter(823)  <=    (tmr_registers(0)(823) and tmr_registers(1)(823)) or                                                             
                            (tmr_registers(1)(823) and tmr_registers(2)(823)) or                                                             
                            (tmr_registers(0)(823) and tmr_registers(2)(823));                                                               
                                                                                                                                         
        local_tmr_voter(824)  <=    (tmr_registers(0)(824) and tmr_registers(1)(824)) or                                                             
                            (tmr_registers(1)(824) and tmr_registers(2)(824)) or                                                             
                            (tmr_registers(0)(824) and tmr_registers(2)(824));                                                               
                                                                                                                                         
        local_tmr_voter(825)  <=    (tmr_registers(0)(825) and tmr_registers(1)(825)) or                                                             
                            (tmr_registers(1)(825) and tmr_registers(2)(825)) or                                                             
                            (tmr_registers(0)(825) and tmr_registers(2)(825));                                                               
                                                                                                                                         
        local_tmr_voter(826)  <=    (tmr_registers(0)(826) and tmr_registers(1)(826)) or                                                             
                            (tmr_registers(1)(826) and tmr_registers(2)(826)) or                                                             
                            (tmr_registers(0)(826) and tmr_registers(2)(826));                                                               
                                                                                                                                         
        local_tmr_voter(827)  <=    (tmr_registers(0)(827) and tmr_registers(1)(827)) or                                                             
                            (tmr_registers(1)(827) and tmr_registers(2)(827)) or                                                             
                            (tmr_registers(0)(827) and tmr_registers(2)(827));                                                               
                                                                                                                                         
        local_tmr_voter(828)  <=    (tmr_registers(0)(828) and tmr_registers(1)(828)) or                                                             
                            (tmr_registers(1)(828) and tmr_registers(2)(828)) or                                                             
                            (tmr_registers(0)(828) and tmr_registers(2)(828));                                                               
                                                                                                                                         
        local_tmr_voter(829)  <=    (tmr_registers(0)(829) and tmr_registers(1)(829)) or                                                             
                            (tmr_registers(1)(829) and tmr_registers(2)(829)) or                                                             
                            (tmr_registers(0)(829) and tmr_registers(2)(829));                                                               
                                                                                                                                         
        local_tmr_voter(830)  <=    (tmr_registers(0)(830) and tmr_registers(1)(830)) or                                                             
                            (tmr_registers(1)(830) and tmr_registers(2)(830)) or                                                             
                            (tmr_registers(0)(830) and tmr_registers(2)(830));                                                               
                                                                                                                                         
        local_tmr_voter(831)  <=    (tmr_registers(0)(831) and tmr_registers(1)(831)) or                                                             
                            (tmr_registers(1)(831) and tmr_registers(2)(831)) or                                                             
                            (tmr_registers(0)(831) and tmr_registers(2)(831));                                                               
                                                                                                                                         
        local_tmr_voter(832)  <=    (tmr_registers(0)(832) and tmr_registers(1)(832)) or                                                             
                            (tmr_registers(1)(832) and tmr_registers(2)(832)) or                                                             
                            (tmr_registers(0)(832) and tmr_registers(2)(832));                                                               
                                                                                                                                         
        local_tmr_voter(833)  <=    (tmr_registers(0)(833) and tmr_registers(1)(833)) or                                                             
                            (tmr_registers(1)(833) and tmr_registers(2)(833)) or                                                             
                            (tmr_registers(0)(833) and tmr_registers(2)(833));                                                               
                                                                                                                                         
        local_tmr_voter(834)  <=    (tmr_registers(0)(834) and tmr_registers(1)(834)) or                                                             
                            (tmr_registers(1)(834) and tmr_registers(2)(834)) or                                                             
                            (tmr_registers(0)(834) and tmr_registers(2)(834));                                                               
                                                                                                                                         
        local_tmr_voter(835)  <=    (tmr_registers(0)(835) and tmr_registers(1)(835)) or                                                             
                            (tmr_registers(1)(835) and tmr_registers(2)(835)) or                                                             
                            (tmr_registers(0)(835) and tmr_registers(2)(835));                                                               
                                                                                                                                         
        local_tmr_voter(836)  <=    (tmr_registers(0)(836) and tmr_registers(1)(836)) or                                                             
                            (tmr_registers(1)(836) and tmr_registers(2)(836)) or                                                             
                            (tmr_registers(0)(836) and tmr_registers(2)(836));                                                               
                                                                                                                                         
        local_tmr_voter(837)  <=    (tmr_registers(0)(837) and tmr_registers(1)(837)) or                                                             
                            (tmr_registers(1)(837) and tmr_registers(2)(837)) or                                                             
                            (tmr_registers(0)(837) and tmr_registers(2)(837));                                                               
                                                                                                                                         
        local_tmr_voter(838)  <=    (tmr_registers(0)(838) and tmr_registers(1)(838)) or                                                             
                            (tmr_registers(1)(838) and tmr_registers(2)(838)) or                                                             
                            (tmr_registers(0)(838) and tmr_registers(2)(838));                                                               
                                                                                                                                         
        local_tmr_voter(839)  <=    (tmr_registers(0)(839) and tmr_registers(1)(839)) or                                                             
                            (tmr_registers(1)(839) and tmr_registers(2)(839)) or                                                             
                            (tmr_registers(0)(839) and tmr_registers(2)(839));                                                               
                                                                                                                                         
        local_tmr_voter(840)  <=    (tmr_registers(0)(840) and tmr_registers(1)(840)) or                                                             
                            (tmr_registers(1)(840) and tmr_registers(2)(840)) or                                                             
                            (tmr_registers(0)(840) and tmr_registers(2)(840));                                                               
                                                                                                                                         
        local_tmr_voter(841)  <=    (tmr_registers(0)(841) and tmr_registers(1)(841)) or                                                             
                            (tmr_registers(1)(841) and tmr_registers(2)(841)) or                                                             
                            (tmr_registers(0)(841) and tmr_registers(2)(841));                                                               
                                                                                                                                         
        local_tmr_voter(842)  <=    (tmr_registers(0)(842) and tmr_registers(1)(842)) or                                                             
                            (tmr_registers(1)(842) and tmr_registers(2)(842)) or                                                             
                            (tmr_registers(0)(842) and tmr_registers(2)(842));                                                               
                                                                                                                                         
        local_tmr_voter(843)  <=    (tmr_registers(0)(843) and tmr_registers(1)(843)) or                                                             
                            (tmr_registers(1)(843) and tmr_registers(2)(843)) or                                                             
                            (tmr_registers(0)(843) and tmr_registers(2)(843));                                                               
                                                                                                                                         
        local_tmr_voter(844)  <=    (tmr_registers(0)(844) and tmr_registers(1)(844)) or                                                             
                            (tmr_registers(1)(844) and tmr_registers(2)(844)) or                                                             
                            (tmr_registers(0)(844) and tmr_registers(2)(844));                                                               
                                                                                                                                         
        local_tmr_voter(845)  <=    (tmr_registers(0)(845) and tmr_registers(1)(845)) or                                                             
                            (tmr_registers(1)(845) and tmr_registers(2)(845)) or                                                             
                            (tmr_registers(0)(845) and tmr_registers(2)(845));                                                               
                                                                                                                                         
        local_tmr_voter(846)  <=    (tmr_registers(0)(846) and tmr_registers(1)(846)) or                                                             
                            (tmr_registers(1)(846) and tmr_registers(2)(846)) or                                                             
                            (tmr_registers(0)(846) and tmr_registers(2)(846));                                                               
                                                                                                                                         
        local_tmr_voter(847)  <=    (tmr_registers(0)(847) and tmr_registers(1)(847)) or                                                             
                            (tmr_registers(1)(847) and tmr_registers(2)(847)) or                                                             
                            (tmr_registers(0)(847) and tmr_registers(2)(847));                                                               
                                                                                                                                         
        local_tmr_voter(848)  <=    (tmr_registers(0)(848) and tmr_registers(1)(848)) or                                                             
                            (tmr_registers(1)(848) and tmr_registers(2)(848)) or                                                             
                            (tmr_registers(0)(848) and tmr_registers(2)(848));                                                               
                                                                                                                                         
        local_tmr_voter(849)  <=    (tmr_registers(0)(849) and tmr_registers(1)(849)) or                                                             
                            (tmr_registers(1)(849) and tmr_registers(2)(849)) or                                                             
                            (tmr_registers(0)(849) and tmr_registers(2)(849));                                                               
                                                                                                                                         
        local_tmr_voter(850)  <=    (tmr_registers(0)(850) and tmr_registers(1)(850)) or                                                             
                            (tmr_registers(1)(850) and tmr_registers(2)(850)) or                                                             
                            (tmr_registers(0)(850) and tmr_registers(2)(850));                                                               
                                                                                                                                         
        local_tmr_voter(851)  <=    (tmr_registers(0)(851) and tmr_registers(1)(851)) or                                                             
                            (tmr_registers(1)(851) and tmr_registers(2)(851)) or                                                             
                            (tmr_registers(0)(851) and tmr_registers(2)(851));                                                               
                                                                                                                                         
        local_tmr_voter(852)  <=    (tmr_registers(0)(852) and tmr_registers(1)(852)) or                                                             
                            (tmr_registers(1)(852) and tmr_registers(2)(852)) or                                                             
                            (tmr_registers(0)(852) and tmr_registers(2)(852));                                                               
                                                                                                                                         
        local_tmr_voter(853)  <=    (tmr_registers(0)(853) and tmr_registers(1)(853)) or                                                             
                            (tmr_registers(1)(853) and tmr_registers(2)(853)) or                                                             
                            (tmr_registers(0)(853) and tmr_registers(2)(853));                                                               
                                                                                                                                         
        local_tmr_voter(854)  <=    (tmr_registers(0)(854) and tmr_registers(1)(854)) or                                                             
                            (tmr_registers(1)(854) and tmr_registers(2)(854)) or                                                             
                            (tmr_registers(0)(854) and tmr_registers(2)(854));                                                               
                                                                                                                                         
        local_tmr_voter(855)  <=    (tmr_registers(0)(855) and tmr_registers(1)(855)) or                                                             
                            (tmr_registers(1)(855) and tmr_registers(2)(855)) or                                                             
                            (tmr_registers(0)(855) and tmr_registers(2)(855));                                                               
                                                                                                                                         
        local_tmr_voter(856)  <=    (tmr_registers(0)(856) and tmr_registers(1)(856)) or                                                             
                            (tmr_registers(1)(856) and tmr_registers(2)(856)) or                                                             
                            (tmr_registers(0)(856) and tmr_registers(2)(856));                                                               
                                                                                                                                         
        local_tmr_voter(857)  <=    (tmr_registers(0)(857) and tmr_registers(1)(857)) or                                                             
                            (tmr_registers(1)(857) and tmr_registers(2)(857)) or                                                             
                            (tmr_registers(0)(857) and tmr_registers(2)(857));                                                               
                                                                                                                                         
        local_tmr_voter(858)  <=    (tmr_registers(0)(858) and tmr_registers(1)(858)) or                                                             
                            (tmr_registers(1)(858) and tmr_registers(2)(858)) or                                                             
                            (tmr_registers(0)(858) and tmr_registers(2)(858));                                                               
                                                                                                                                         
        local_tmr_voter(859)  <=    (tmr_registers(0)(859) and tmr_registers(1)(859)) or                                                             
                            (tmr_registers(1)(859) and tmr_registers(2)(859)) or                                                             
                            (tmr_registers(0)(859) and tmr_registers(2)(859));                                                               
                                                                                                                                         
        local_tmr_voter(860)  <=    (tmr_registers(0)(860) and tmr_registers(1)(860)) or                                                             
                            (tmr_registers(1)(860) and tmr_registers(2)(860)) or                                                             
                            (tmr_registers(0)(860) and tmr_registers(2)(860));                                                               
                                                                                                                                         
        local_tmr_voter(861)  <=    (tmr_registers(0)(861) and tmr_registers(1)(861)) or                                                             
                            (tmr_registers(1)(861) and tmr_registers(2)(861)) or                                                             
                            (tmr_registers(0)(861) and tmr_registers(2)(861));                                                               
                                                                                                                                         
        local_tmr_voter(862)  <=    (tmr_registers(0)(862) and tmr_registers(1)(862)) or                                                             
                            (tmr_registers(1)(862) and tmr_registers(2)(862)) or                                                             
                            (tmr_registers(0)(862) and tmr_registers(2)(862));                                                               
                                                                                                                                         
        local_tmr_voter(863)  <=    (tmr_registers(0)(863) and tmr_registers(1)(863)) or                                                             
                            (tmr_registers(1)(863) and tmr_registers(2)(863)) or                                                             
                            (tmr_registers(0)(863) and tmr_registers(2)(863));                                                               
                                                                                                                                         
        local_tmr_voter(864)  <=    (tmr_registers(0)(864) and tmr_registers(1)(864)) or                                                             
                            (tmr_registers(1)(864) and tmr_registers(2)(864)) or                                                             
                            (tmr_registers(0)(864) and tmr_registers(2)(864));                                                               
                                                                                                                                         
        local_tmr_voter(865)  <=    (tmr_registers(0)(865) and tmr_registers(1)(865)) or                                                             
                            (tmr_registers(1)(865) and tmr_registers(2)(865)) or                                                             
                            (tmr_registers(0)(865) and tmr_registers(2)(865));                                                               
                                                                                                                                         
        local_tmr_voter(866)  <=    (tmr_registers(0)(866) and tmr_registers(1)(866)) or                                                             
                            (tmr_registers(1)(866) and tmr_registers(2)(866)) or                                                             
                            (tmr_registers(0)(866) and tmr_registers(2)(866));                                                               
                                                                                                                                         
        local_tmr_voter(867)  <=    (tmr_registers(0)(867) and tmr_registers(1)(867)) or                                                             
                            (tmr_registers(1)(867) and tmr_registers(2)(867)) or                                                             
                            (tmr_registers(0)(867) and tmr_registers(2)(867));                                                               
                                                                                                                                         
        local_tmr_voter(868)  <=    (tmr_registers(0)(868) and tmr_registers(1)(868)) or                                                             
                            (tmr_registers(1)(868) and tmr_registers(2)(868)) or                                                             
                            (tmr_registers(0)(868) and tmr_registers(2)(868));                                                               
                                                                                                                                         
        local_tmr_voter(869)  <=    (tmr_registers(0)(869) and tmr_registers(1)(869)) or                                                             
                            (tmr_registers(1)(869) and tmr_registers(2)(869)) or                                                             
                            (tmr_registers(0)(869) and tmr_registers(2)(869));                                                               
                                                                                                                                         
        local_tmr_voter(870)  <=    (tmr_registers(0)(870) and tmr_registers(1)(870)) or                                                             
                            (tmr_registers(1)(870) and tmr_registers(2)(870)) or                                                             
                            (tmr_registers(0)(870) and tmr_registers(2)(870));                                                               
                                                                                                                                         
        local_tmr_voter(871)  <=    (tmr_registers(0)(871) and tmr_registers(1)(871)) or                                                             
                            (tmr_registers(1)(871) and tmr_registers(2)(871)) or                                                             
                            (tmr_registers(0)(871) and tmr_registers(2)(871));                                                               
                                                                                                                                         
        local_tmr_voter(872)  <=    (tmr_registers(0)(872) and tmr_registers(1)(872)) or                                                             
                            (tmr_registers(1)(872) and tmr_registers(2)(872)) or                                                             
                            (tmr_registers(0)(872) and tmr_registers(2)(872));                                                               
                                                                                                                                         
        local_tmr_voter(873)  <=    (tmr_registers(0)(873) and tmr_registers(1)(873)) or                                                             
                            (tmr_registers(1)(873) and tmr_registers(2)(873)) or                                                             
                            (tmr_registers(0)(873) and tmr_registers(2)(873));                                                               
                                                                                                                                         
        local_tmr_voter(874)  <=    (tmr_registers(0)(874) and tmr_registers(1)(874)) or                                                             
                            (tmr_registers(1)(874) and tmr_registers(2)(874)) or                                                             
                            (tmr_registers(0)(874) and tmr_registers(2)(874));                                                               
                                                                                                                                         
        local_tmr_voter(875)  <=    (tmr_registers(0)(875) and tmr_registers(1)(875)) or                                                             
                            (tmr_registers(1)(875) and tmr_registers(2)(875)) or                                                             
                            (tmr_registers(0)(875) and tmr_registers(2)(875));                                                               
                                                                                                                                         
        local_tmr_voter(876)  <=    (tmr_registers(0)(876) and tmr_registers(1)(876)) or                                                             
                            (tmr_registers(1)(876) and tmr_registers(2)(876)) or                                                             
                            (tmr_registers(0)(876) and tmr_registers(2)(876));                                                               
                                                                                                                                         
        local_tmr_voter(877)  <=    (tmr_registers(0)(877) and tmr_registers(1)(877)) or                                                             
                            (tmr_registers(1)(877) and tmr_registers(2)(877)) or                                                             
                            (tmr_registers(0)(877) and tmr_registers(2)(877));                                                               
                                                                                                                                         
        local_tmr_voter(878)  <=    (tmr_registers(0)(878) and tmr_registers(1)(878)) or                                                             
                            (tmr_registers(1)(878) and tmr_registers(2)(878)) or                                                             
                            (tmr_registers(0)(878) and tmr_registers(2)(878));                                                               
                                                                                                                                         
        local_tmr_voter(879)  <=    (tmr_registers(0)(879) and tmr_registers(1)(879)) or                                                             
                            (tmr_registers(1)(879) and tmr_registers(2)(879)) or                                                             
                            (tmr_registers(0)(879) and tmr_registers(2)(879));                                                               
                                                                                                                                         
        local_tmr_voter(880)  <=    (tmr_registers(0)(880) and tmr_registers(1)(880)) or                                                             
                            (tmr_registers(1)(880) and tmr_registers(2)(880)) or                                                             
                            (tmr_registers(0)(880) and tmr_registers(2)(880));                                                               
                                                                                                                                         
        local_tmr_voter(881)  <=    (tmr_registers(0)(881) and tmr_registers(1)(881)) or                                                             
                            (tmr_registers(1)(881) and tmr_registers(2)(881)) or                                                             
                            (tmr_registers(0)(881) and tmr_registers(2)(881));                                                               
                                                                                                                                         
        local_tmr_voter(882)  <=    (tmr_registers(0)(882) and tmr_registers(1)(882)) or                                                             
                            (tmr_registers(1)(882) and tmr_registers(2)(882)) or                                                             
                            (tmr_registers(0)(882) and tmr_registers(2)(882));                                                               
                                                                                                                                         
        local_tmr_voter(883)  <=    (tmr_registers(0)(883) and tmr_registers(1)(883)) or                                                             
                            (tmr_registers(1)(883) and tmr_registers(2)(883)) or                                                             
                            (tmr_registers(0)(883) and tmr_registers(2)(883));                                                               
                                                                                                                                         
        local_tmr_voter(884)  <=    (tmr_registers(0)(884) and tmr_registers(1)(884)) or                                                             
                            (tmr_registers(1)(884) and tmr_registers(2)(884)) or                                                             
                            (tmr_registers(0)(884) and tmr_registers(2)(884));                                                               
                                                                                                                                         
        local_tmr_voter(885)  <=    (tmr_registers(0)(885) and tmr_registers(1)(885)) or                                                             
                            (tmr_registers(1)(885) and tmr_registers(2)(885)) or                                                             
                            (tmr_registers(0)(885) and tmr_registers(2)(885));                                                               
                                                                                                                                         
        local_tmr_voter(886)  <=    (tmr_registers(0)(886) and tmr_registers(1)(886)) or                                                             
                            (tmr_registers(1)(886) and tmr_registers(2)(886)) or                                                             
                            (tmr_registers(0)(886) and tmr_registers(2)(886));                                                               
                                                                                                                                         
        local_tmr_voter(887)  <=    (tmr_registers(0)(887) and tmr_registers(1)(887)) or                                                             
                            (tmr_registers(1)(887) and tmr_registers(2)(887)) or                                                             
                            (tmr_registers(0)(887) and tmr_registers(2)(887));                                                               
                                                                                                                                         
        local_tmr_voter(888)  <=    (tmr_registers(0)(888) and tmr_registers(1)(888)) or                                                             
                            (tmr_registers(1)(888) and tmr_registers(2)(888)) or                                                             
                            (tmr_registers(0)(888) and tmr_registers(2)(888));                                                               
                                                                                                                                         
        local_tmr_voter(889)  <=    (tmr_registers(0)(889) and tmr_registers(1)(889)) or                                                             
                            (tmr_registers(1)(889) and tmr_registers(2)(889)) or                                                             
                            (tmr_registers(0)(889) and tmr_registers(2)(889));                                                               
                                                                                                                                         
        local_tmr_voter(890)  <=    (tmr_registers(0)(890) and tmr_registers(1)(890)) or                                                             
                            (tmr_registers(1)(890) and tmr_registers(2)(890)) or                                                             
                            (tmr_registers(0)(890) and tmr_registers(2)(890));                                                               
                                                                                                                                         
        local_tmr_voter(891)  <=    (tmr_registers(0)(891) and tmr_registers(1)(891)) or                                                             
                            (tmr_registers(1)(891) and tmr_registers(2)(891)) or                                                             
                            (tmr_registers(0)(891) and tmr_registers(2)(891));                                                               
                                                                                                                                         
        local_tmr_voter(892)  <=    (tmr_registers(0)(892) and tmr_registers(1)(892)) or                                                             
                            (tmr_registers(1)(892) and tmr_registers(2)(892)) or                                                             
                            (tmr_registers(0)(892) and tmr_registers(2)(892));                                                               
                                                                                                                                         
        local_tmr_voter(893)  <=    (tmr_registers(0)(893) and tmr_registers(1)(893)) or                                                             
                            (tmr_registers(1)(893) and tmr_registers(2)(893)) or                                                             
                            (tmr_registers(0)(893) and tmr_registers(2)(893));                                                               
                                                                                                                                         
        local_tmr_voter(894)  <=    (tmr_registers(0)(894) and tmr_registers(1)(894)) or                                                             
                            (tmr_registers(1)(894) and tmr_registers(2)(894)) or                                                             
                            (tmr_registers(0)(894) and tmr_registers(2)(894));                                                               
                                                                                                                                         
        local_tmr_voter(895)  <=    (tmr_registers(0)(895) and tmr_registers(1)(895)) or                                                             
                            (tmr_registers(1)(895) and tmr_registers(2)(895)) or                                                             
                            (tmr_registers(0)(895) and tmr_registers(2)(895));                                                               
                                                                                                                                         
        local_tmr_voter(896)  <=    (tmr_registers(0)(896) and tmr_registers(1)(896)) or                                                             
                            (tmr_registers(1)(896) and tmr_registers(2)(896)) or                                                             
                            (tmr_registers(0)(896) and tmr_registers(2)(896));                                                               
                                                                                                                                         
        local_tmr_voter(897)  <=    (tmr_registers(0)(897) and tmr_registers(1)(897)) or                                                             
                            (tmr_registers(1)(897) and tmr_registers(2)(897)) or                                                             
                            (tmr_registers(0)(897) and tmr_registers(2)(897));                                                               
                                                                                                                                         
        local_tmr_voter(898)  <=    (tmr_registers(0)(898) and tmr_registers(1)(898)) or                                                             
                            (tmr_registers(1)(898) and tmr_registers(2)(898)) or                                                             
                            (tmr_registers(0)(898) and tmr_registers(2)(898));                                                               
                                                                                                                                         
        local_tmr_voter(899)  <=    (tmr_registers(0)(899) and tmr_registers(1)(899)) or                                                             
                            (tmr_registers(1)(899) and tmr_registers(2)(899)) or                                                             
                            (tmr_registers(0)(899) and tmr_registers(2)(899));                                                               
                                                                                                                                         
        local_tmr_voter(900)  <=    (tmr_registers(0)(900) and tmr_registers(1)(900)) or                                                             
                            (tmr_registers(1)(900) and tmr_registers(2)(900)) or                                                             
                            (tmr_registers(0)(900) and tmr_registers(2)(900));                                                               
                                                                                                                                         
        local_tmr_voter(901)  <=    (tmr_registers(0)(901) and tmr_registers(1)(901)) or                                                             
                            (tmr_registers(1)(901) and tmr_registers(2)(901)) or                                                             
                            (tmr_registers(0)(901) and tmr_registers(2)(901));                                                               
                                                                                                                                         
        local_tmr_voter(902)  <=    (tmr_registers(0)(902) and tmr_registers(1)(902)) or                                                             
                            (tmr_registers(1)(902) and tmr_registers(2)(902)) or                                                             
                            (tmr_registers(0)(902) and tmr_registers(2)(902));                                                               
                                                                                                                                         
        local_tmr_voter(903)  <=    (tmr_registers(0)(903) and tmr_registers(1)(903)) or                                                             
                            (tmr_registers(1)(903) and tmr_registers(2)(903)) or                                                             
                            (tmr_registers(0)(903) and tmr_registers(2)(903));                                                               
                                                                                                                                         
        local_tmr_voter(904)  <=    (tmr_registers(0)(904) and tmr_registers(1)(904)) or                                                             
                            (tmr_registers(1)(904) and tmr_registers(2)(904)) or                                                             
                            (tmr_registers(0)(904) and tmr_registers(2)(904));                                                               
                                                                                                                                         
        local_tmr_voter(905)  <=    (tmr_registers(0)(905) and tmr_registers(1)(905)) or                                                             
                            (tmr_registers(1)(905) and tmr_registers(2)(905)) or                                                             
                            (tmr_registers(0)(905) and tmr_registers(2)(905));                                                               
                                                                                                                                         
        local_tmr_voter(906)  <=    (tmr_registers(0)(906) and tmr_registers(1)(906)) or                                                             
                            (tmr_registers(1)(906) and tmr_registers(2)(906)) or                                                             
                            (tmr_registers(0)(906) and tmr_registers(2)(906));                                                               
                                                                                                                                         
        local_tmr_voter(907)  <=    (tmr_registers(0)(907) and tmr_registers(1)(907)) or                                                             
                            (tmr_registers(1)(907) and tmr_registers(2)(907)) or                                                             
                            (tmr_registers(0)(907) and tmr_registers(2)(907));                                                               
                                                                                                                                         
        local_tmr_voter(908)  <=    (tmr_registers(0)(908) and tmr_registers(1)(908)) or                                                             
                            (tmr_registers(1)(908) and tmr_registers(2)(908)) or                                                             
                            (tmr_registers(0)(908) and tmr_registers(2)(908));                                                               
                                                                                                                                         
        local_tmr_voter(909)  <=    (tmr_registers(0)(909) and tmr_registers(1)(909)) or                                                             
                            (tmr_registers(1)(909) and tmr_registers(2)(909)) or                                                             
                            (tmr_registers(0)(909) and tmr_registers(2)(909));                                                               
                                                                                                                                         
        local_tmr_voter(910)  <=    (tmr_registers(0)(910) and tmr_registers(1)(910)) or                                                             
                            (tmr_registers(1)(910) and tmr_registers(2)(910)) or                                                             
                            (tmr_registers(0)(910) and tmr_registers(2)(910));                                                               
                                                                                                                                         
        local_tmr_voter(911)  <=    (tmr_registers(0)(911) and tmr_registers(1)(911)) or                                                             
                            (tmr_registers(1)(911) and tmr_registers(2)(911)) or                                                             
                            (tmr_registers(0)(911) and tmr_registers(2)(911));                                                               
                                                                                                                                         
        local_tmr_voter(912)  <=    (tmr_registers(0)(912) and tmr_registers(1)(912)) or                                                             
                            (tmr_registers(1)(912) and tmr_registers(2)(912)) or                                                             
                            (tmr_registers(0)(912) and tmr_registers(2)(912));                                                               
                                                                                                                                         
        local_tmr_voter(913)  <=    (tmr_registers(0)(913) and tmr_registers(1)(913)) or                                                             
                            (tmr_registers(1)(913) and tmr_registers(2)(913)) or                                                             
                            (tmr_registers(0)(913) and tmr_registers(2)(913));                                                               
                                                                                                                                         
        local_tmr_voter(914)  <=    (tmr_registers(0)(914) and tmr_registers(1)(914)) or                                                             
                            (tmr_registers(1)(914) and tmr_registers(2)(914)) or                                                             
                            (tmr_registers(0)(914) and tmr_registers(2)(914));                                                               
                                                                                                                                         
        local_tmr_voter(915)  <=    (tmr_registers(0)(915) and tmr_registers(1)(915)) or                                                             
                            (tmr_registers(1)(915) and tmr_registers(2)(915)) or                                                             
                            (tmr_registers(0)(915) and tmr_registers(2)(915));                                                               
                                                                                                                                         
        local_tmr_voter(916)  <=    (tmr_registers(0)(916) and tmr_registers(1)(916)) or                                                             
                            (tmr_registers(1)(916) and tmr_registers(2)(916)) or                                                             
                            (tmr_registers(0)(916) and tmr_registers(2)(916));                                                               
                                                                                                                                         
        local_tmr_voter(917)  <=    (tmr_registers(0)(917) and tmr_registers(1)(917)) or                                                             
                            (tmr_registers(1)(917) and tmr_registers(2)(917)) or                                                             
                            (tmr_registers(0)(917) and tmr_registers(2)(917));                                                               
                                                                                                                                         
        local_tmr_voter(918)  <=    (tmr_registers(0)(918) and tmr_registers(1)(918)) or                                                             
                            (tmr_registers(1)(918) and tmr_registers(2)(918)) or                                                             
                            (tmr_registers(0)(918) and tmr_registers(2)(918));                                                               
                                                                                                                                         
        local_tmr_voter(919)  <=    (tmr_registers(0)(919) and tmr_registers(1)(919)) or                                                             
                            (tmr_registers(1)(919) and tmr_registers(2)(919)) or                                                             
                            (tmr_registers(0)(919) and tmr_registers(2)(919));                                                               
                                                                                                                                         
        local_tmr_voter(920)  <=    (tmr_registers(0)(920) and tmr_registers(1)(920)) or                                                             
                            (tmr_registers(1)(920) and tmr_registers(2)(920)) or                                                             
                            (tmr_registers(0)(920) and tmr_registers(2)(920));                                                               
                                                                                                                                         
        local_tmr_voter(921)  <=    (tmr_registers(0)(921) and tmr_registers(1)(921)) or                                                             
                            (tmr_registers(1)(921) and tmr_registers(2)(921)) or                                                             
                            (tmr_registers(0)(921) and tmr_registers(2)(921));                                                               
                                                                                                                                         
        local_tmr_voter(922)  <=    (tmr_registers(0)(922) and tmr_registers(1)(922)) or                                                             
                            (tmr_registers(1)(922) and tmr_registers(2)(922)) or                                                             
                            (tmr_registers(0)(922) and tmr_registers(2)(922));                                                               
                                                                                                                                         
        local_tmr_voter(923)  <=    (tmr_registers(0)(923) and tmr_registers(1)(923)) or                                                             
                            (tmr_registers(1)(923) and tmr_registers(2)(923)) or                                                             
                            (tmr_registers(0)(923) and tmr_registers(2)(923));                                                               
                                                                                                                                         
        local_tmr_voter(924)  <=    (tmr_registers(0)(924) and tmr_registers(1)(924)) or                                                             
                            (tmr_registers(1)(924) and tmr_registers(2)(924)) or                                                             
                            (tmr_registers(0)(924) and tmr_registers(2)(924));                                                               
                                                                                                                                         
        local_tmr_voter(925)  <=    (tmr_registers(0)(925) and tmr_registers(1)(925)) or                                                             
                            (tmr_registers(1)(925) and tmr_registers(2)(925)) or                                                             
                            (tmr_registers(0)(925) and tmr_registers(2)(925));                                                               
                                                                                                                                         
        local_tmr_voter(926)  <=    (tmr_registers(0)(926) and tmr_registers(1)(926)) or                                                             
                            (tmr_registers(1)(926) and tmr_registers(2)(926)) or                                                             
                            (tmr_registers(0)(926) and tmr_registers(2)(926));                                                               
                                                                                                                                         
        local_tmr_voter(927)  <=    (tmr_registers(0)(927) and tmr_registers(1)(927)) or                                                             
                            (tmr_registers(1)(927) and tmr_registers(2)(927)) or                                                             
                            (tmr_registers(0)(927) and tmr_registers(2)(927));                                                               
                                                                                                                                         
        local_tmr_voter(928)  <=    (tmr_registers(0)(928) and tmr_registers(1)(928)) or                                                             
                            (tmr_registers(1)(928) and tmr_registers(2)(928)) or                                                             
                            (tmr_registers(0)(928) and tmr_registers(2)(928));                                                               
                                                                                                                                         
        local_tmr_voter(929)  <=    (tmr_registers(0)(929) and tmr_registers(1)(929)) or                                                             
                            (tmr_registers(1)(929) and tmr_registers(2)(929)) or                                                             
                            (tmr_registers(0)(929) and tmr_registers(2)(929));                                                               
                                                                                                                                         
        local_tmr_voter(930)  <=    (tmr_registers(0)(930) and tmr_registers(1)(930)) or                                                             
                            (tmr_registers(1)(930) and tmr_registers(2)(930)) or                                                             
                            (tmr_registers(0)(930) and tmr_registers(2)(930));                                                               
                                                                                                                                         
        local_tmr_voter(931)  <=    (tmr_registers(0)(931) and tmr_registers(1)(931)) or                                                             
                            (tmr_registers(1)(931) and tmr_registers(2)(931)) or                                                             
                            (tmr_registers(0)(931) and tmr_registers(2)(931));                                                               
                                                                                                                                         
        local_tmr_voter(932)  <=    (tmr_registers(0)(932) and tmr_registers(1)(932)) or                                                             
                            (tmr_registers(1)(932) and tmr_registers(2)(932)) or                                                             
                            (tmr_registers(0)(932) and tmr_registers(2)(932));                                                               
                                                                                                                                         
        local_tmr_voter(933)  <=    (tmr_registers(0)(933) and tmr_registers(1)(933)) or                                                             
                            (tmr_registers(1)(933) and tmr_registers(2)(933)) or                                                             
                            (tmr_registers(0)(933) and tmr_registers(2)(933));                                                               
                                                                                                                                         
        local_tmr_voter(934)  <=    (tmr_registers(0)(934) and tmr_registers(1)(934)) or                                                             
                            (tmr_registers(1)(934) and tmr_registers(2)(934)) or                                                             
                            (tmr_registers(0)(934) and tmr_registers(2)(934));                                                               
                                                                                                                                         
        local_tmr_voter(935)  <=    (tmr_registers(0)(935) and tmr_registers(1)(935)) or                                                             
                            (tmr_registers(1)(935) and tmr_registers(2)(935)) or                                                             
                            (tmr_registers(0)(935) and tmr_registers(2)(935));                                                               
                                                                                                                                         
        local_tmr_voter(936)  <=    (tmr_registers(0)(936) and tmr_registers(1)(936)) or                                                             
                            (tmr_registers(1)(936) and tmr_registers(2)(936)) or                                                             
                            (tmr_registers(0)(936) and tmr_registers(2)(936));                                                               
                                                                                                                                         
        local_tmr_voter(937)  <=    (tmr_registers(0)(937) and tmr_registers(1)(937)) or                                                             
                            (tmr_registers(1)(937) and tmr_registers(2)(937)) or                                                             
                            (tmr_registers(0)(937) and tmr_registers(2)(937));                                                               
                                                                                                                                         
        local_tmr_voter(938)  <=    (tmr_registers(0)(938) and tmr_registers(1)(938)) or                                                             
                            (tmr_registers(1)(938) and tmr_registers(2)(938)) or                                                             
                            (tmr_registers(0)(938) and tmr_registers(2)(938));                                                               
                                                                                                                                         
        local_tmr_voter(939)  <=    (tmr_registers(0)(939) and tmr_registers(1)(939)) or                                                             
                            (tmr_registers(1)(939) and tmr_registers(2)(939)) or                                                             
                            (tmr_registers(0)(939) and tmr_registers(2)(939));                                                               
                                                                                                                                         
        local_tmr_voter(940)  <=    (tmr_registers(0)(940) and tmr_registers(1)(940)) or                                                             
                            (tmr_registers(1)(940) and tmr_registers(2)(940)) or                                                             
                            (tmr_registers(0)(940) and tmr_registers(2)(940));                                                               
                                                                                                                                         
        local_tmr_voter(941)  <=    (tmr_registers(0)(941) and tmr_registers(1)(941)) or                                                             
                            (tmr_registers(1)(941) and tmr_registers(2)(941)) or                                                             
                            (tmr_registers(0)(941) and tmr_registers(2)(941));                                                               
                                                                                                                                         
        local_tmr_voter(942)  <=    (tmr_registers(0)(942) and tmr_registers(1)(942)) or                                                             
                            (tmr_registers(1)(942) and tmr_registers(2)(942)) or                                                             
                            (tmr_registers(0)(942) and tmr_registers(2)(942));                                                               
                                                                                                                                         
        local_tmr_voter(943)  <=    (tmr_registers(0)(943) and tmr_registers(1)(943)) or                                                             
                            (tmr_registers(1)(943) and tmr_registers(2)(943)) or                                                             
                            (tmr_registers(0)(943) and tmr_registers(2)(943));                                                               
                                                                                                                                         
        local_tmr_voter(944)  <=    (tmr_registers(0)(944) and tmr_registers(1)(944)) or                                                             
                            (tmr_registers(1)(944) and tmr_registers(2)(944)) or                                                             
                            (tmr_registers(0)(944) and tmr_registers(2)(944));                                                               
                                                                                                                                         
        local_tmr_voter(945)  <=    (tmr_registers(0)(945) and tmr_registers(1)(945)) or                                                             
                            (tmr_registers(1)(945) and tmr_registers(2)(945)) or                                                             
                            (tmr_registers(0)(945) and tmr_registers(2)(945));                                                               
                                                                                                                                         
        local_tmr_voter(946)  <=    (tmr_registers(0)(946) and tmr_registers(1)(946)) or                                                             
                            (tmr_registers(1)(946) and tmr_registers(2)(946)) or                                                             
                            (tmr_registers(0)(946) and tmr_registers(2)(946));                                                               
                                                                                                                                         
        local_tmr_voter(947)  <=    (tmr_registers(0)(947) and tmr_registers(1)(947)) or                                                             
                            (tmr_registers(1)(947) and tmr_registers(2)(947)) or                                                             
                            (tmr_registers(0)(947) and tmr_registers(2)(947));                                                               
                                                                                                                                         
        local_tmr_voter(948)  <=    (tmr_registers(0)(948) and tmr_registers(1)(948)) or                                                             
                            (tmr_registers(1)(948) and tmr_registers(2)(948)) or                                                             
                            (tmr_registers(0)(948) and tmr_registers(2)(948));                                                               
                                                                                                                                         
        local_tmr_voter(949)  <=    (tmr_registers(0)(949) and tmr_registers(1)(949)) or                                                             
                            (tmr_registers(1)(949) and tmr_registers(2)(949)) or                                                             
                            (tmr_registers(0)(949) and tmr_registers(2)(949));                                                               
                                                                                                                                         
        local_tmr_voter(950)  <=    (tmr_registers(0)(950) and tmr_registers(1)(950)) or                                                             
                            (tmr_registers(1)(950) and tmr_registers(2)(950)) or                                                             
                            (tmr_registers(0)(950) and tmr_registers(2)(950));                                                               
                                                                                                                                         
        local_tmr_voter(951)  <=    (tmr_registers(0)(951) and tmr_registers(1)(951)) or                                                             
                            (tmr_registers(1)(951) and tmr_registers(2)(951)) or                                                             
                            (tmr_registers(0)(951) and tmr_registers(2)(951));                                                               
                                                                                                                                         
        local_tmr_voter(952)  <=    (tmr_registers(0)(952) and tmr_registers(1)(952)) or                                                             
                            (tmr_registers(1)(952) and tmr_registers(2)(952)) or                                                             
                            (tmr_registers(0)(952) and tmr_registers(2)(952));                                                               
                                                                                                                                         
        local_tmr_voter(953)  <=    (tmr_registers(0)(953) and tmr_registers(1)(953)) or                                                             
                            (tmr_registers(1)(953) and tmr_registers(2)(953)) or                                                             
                            (tmr_registers(0)(953) and tmr_registers(2)(953));                                                               
                                                                                                                                         
        local_tmr_voter(954)  <=    (tmr_registers(0)(954) and tmr_registers(1)(954)) or                                                             
                            (tmr_registers(1)(954) and tmr_registers(2)(954)) or                                                             
                            (tmr_registers(0)(954) and tmr_registers(2)(954));                                                               
                                                                                                                                         
        local_tmr_voter(955)  <=    (tmr_registers(0)(955) and tmr_registers(1)(955)) or                                                             
                            (tmr_registers(1)(955) and tmr_registers(2)(955)) or                                                             
                            (tmr_registers(0)(955) and tmr_registers(2)(955));                                                               
                                                                                                                                         
        local_tmr_voter(956)  <=    (tmr_registers(0)(956) and tmr_registers(1)(956)) or                                                             
                            (tmr_registers(1)(956) and tmr_registers(2)(956)) or                                                             
                            (tmr_registers(0)(956) and tmr_registers(2)(956));                                                               
                                                                                                                                         
        local_tmr_voter(957)  <=    (tmr_registers(0)(957) and tmr_registers(1)(957)) or                                                             
                            (tmr_registers(1)(957) and tmr_registers(2)(957)) or                                                             
                            (tmr_registers(0)(957) and tmr_registers(2)(957));                                                               
                                                                                                                                         
        local_tmr_voter(958)  <=    (tmr_registers(0)(958) and tmr_registers(1)(958)) or                                                             
                            (tmr_registers(1)(958) and tmr_registers(2)(958)) or                                                             
                            (tmr_registers(0)(958) and tmr_registers(2)(958));                                                               
                                                                                                                                         
        local_tmr_voter(959)  <=    (tmr_registers(0)(959) and tmr_registers(1)(959)) or                                                             
                            (tmr_registers(1)(959) and tmr_registers(2)(959)) or                                                             
                            (tmr_registers(0)(959) and tmr_registers(2)(959));                                                               
                                                                                                                                         
        local_tmr_voter(960)  <=    (tmr_registers(0)(960) and tmr_registers(1)(960)) or                                                             
                            (tmr_registers(1)(960) and tmr_registers(2)(960)) or                                                             
                            (tmr_registers(0)(960) and tmr_registers(2)(960));                                                               
                                                                                                                                         
        local_tmr_voter(961)  <=    (tmr_registers(0)(961) and tmr_registers(1)(961)) or                                                             
                            (tmr_registers(1)(961) and tmr_registers(2)(961)) or                                                             
                            (tmr_registers(0)(961) and tmr_registers(2)(961));                                                               
                                                                                                                                         
        local_tmr_voter(962)  <=    (tmr_registers(0)(962) and tmr_registers(1)(962)) or                                                             
                            (tmr_registers(1)(962) and tmr_registers(2)(962)) or                                                             
                            (tmr_registers(0)(962) and tmr_registers(2)(962));                                                               
                                                                                                                                         
        local_tmr_voter(963)  <=    (tmr_registers(0)(963) and tmr_registers(1)(963)) or                                                             
                            (tmr_registers(1)(963) and tmr_registers(2)(963)) or                                                             
                            (tmr_registers(0)(963) and tmr_registers(2)(963));                                                               
                                                                                                                                         
        local_tmr_voter(964)  <=    (tmr_registers(0)(964) and tmr_registers(1)(964)) or                                                             
                            (tmr_registers(1)(964) and tmr_registers(2)(964)) or                                                             
                            (tmr_registers(0)(964) and tmr_registers(2)(964));                                                               
                                                                                                                                         
        local_tmr_voter(965)  <=    (tmr_registers(0)(965) and tmr_registers(1)(965)) or                                                             
                            (tmr_registers(1)(965) and tmr_registers(2)(965)) or                                                             
                            (tmr_registers(0)(965) and tmr_registers(2)(965));                                                               
                                                                                                                                         
        local_tmr_voter(966)  <=    (tmr_registers(0)(966) and tmr_registers(1)(966)) or                                                             
                            (tmr_registers(1)(966) and tmr_registers(2)(966)) or                                                             
                            (tmr_registers(0)(966) and tmr_registers(2)(966));                                                               
                                                                                                                                         
        local_tmr_voter(967)  <=    (tmr_registers(0)(967) and tmr_registers(1)(967)) or                                                             
                            (tmr_registers(1)(967) and tmr_registers(2)(967)) or                                                             
                            (tmr_registers(0)(967) and tmr_registers(2)(967));                                                               
                                                                                                                                         
        local_tmr_voter(968)  <=    (tmr_registers(0)(968) and tmr_registers(1)(968)) or                                                             
                            (tmr_registers(1)(968) and tmr_registers(2)(968)) or                                                             
                            (tmr_registers(0)(968) and tmr_registers(2)(968));                                                               
                                                                                                                                         
        local_tmr_voter(969)  <=    (tmr_registers(0)(969) and tmr_registers(1)(969)) or                                                             
                            (tmr_registers(1)(969) and tmr_registers(2)(969)) or                                                             
                            (tmr_registers(0)(969) and tmr_registers(2)(969));                                                               
                                                                                                                                         
        local_tmr_voter(970)  <=    (tmr_registers(0)(970) and tmr_registers(1)(970)) or                                                             
                            (tmr_registers(1)(970) and tmr_registers(2)(970)) or                                                             
                            (tmr_registers(0)(970) and tmr_registers(2)(970));                                                               
                                                                                                                                         
        local_tmr_voter(971)  <=    (tmr_registers(0)(971) and tmr_registers(1)(971)) or                                                             
                            (tmr_registers(1)(971) and tmr_registers(2)(971)) or                                                             
                            (tmr_registers(0)(971) and tmr_registers(2)(971));                                                               
                                                                                                                                         
        local_tmr_voter(972)  <=    (tmr_registers(0)(972) and tmr_registers(1)(972)) or                                                             
                            (tmr_registers(1)(972) and tmr_registers(2)(972)) or                                                             
                            (tmr_registers(0)(972) and tmr_registers(2)(972));                                                               
                                                                                                                                         
        local_tmr_voter(973)  <=    (tmr_registers(0)(973) and tmr_registers(1)(973)) or                                                             
                            (tmr_registers(1)(973) and tmr_registers(2)(973)) or                                                             
                            (tmr_registers(0)(973) and tmr_registers(2)(973));                                                               
                                                                                                                                         
        local_tmr_voter(974)  <=    (tmr_registers(0)(974) and tmr_registers(1)(974)) or                                                             
                            (tmr_registers(1)(974) and tmr_registers(2)(974)) or                                                             
                            (tmr_registers(0)(974) and tmr_registers(2)(974));                                                               
                                                                                                                                         
        local_tmr_voter(975)  <=    (tmr_registers(0)(975) and tmr_registers(1)(975)) or                                                             
                            (tmr_registers(1)(975) and tmr_registers(2)(975)) or                                                             
                            (tmr_registers(0)(975) and tmr_registers(2)(975));                                                               
                                                                                                                                         
        local_tmr_voter(976)  <=    (tmr_registers(0)(976) and tmr_registers(1)(976)) or                                                             
                            (tmr_registers(1)(976) and tmr_registers(2)(976)) or                                                             
                            (tmr_registers(0)(976) and tmr_registers(2)(976));                                                               
                                                                                                                                         
        local_tmr_voter(977)  <=    (tmr_registers(0)(977) and tmr_registers(1)(977)) or                                                             
                            (tmr_registers(1)(977) and tmr_registers(2)(977)) or                                                             
                            (tmr_registers(0)(977) and tmr_registers(2)(977));                                                               
                                                                                                                                         
        local_tmr_voter(978)  <=    (tmr_registers(0)(978) and tmr_registers(1)(978)) or                                                             
                            (tmr_registers(1)(978) and tmr_registers(2)(978)) or                                                             
                            (tmr_registers(0)(978) and tmr_registers(2)(978));                                                               
                                                                                                                                         
        local_tmr_voter(979)  <=    (tmr_registers(0)(979) and tmr_registers(1)(979)) or                                                             
                            (tmr_registers(1)(979) and tmr_registers(2)(979)) or                                                             
                            (tmr_registers(0)(979) and tmr_registers(2)(979));                                                               
                                                                                                                                         
        local_tmr_voter(980)  <=    (tmr_registers(0)(980) and tmr_registers(1)(980)) or                                                             
                            (tmr_registers(1)(980) and tmr_registers(2)(980)) or                                                             
                            (tmr_registers(0)(980) and tmr_registers(2)(980));                                                               
                                                                                                                                         
        local_tmr_voter(981)  <=    (tmr_registers(0)(981) and tmr_registers(1)(981)) or                                                             
                            (tmr_registers(1)(981) and tmr_registers(2)(981)) or                                                             
                            (tmr_registers(0)(981) and tmr_registers(2)(981));                                                               
                                                                                                                                         
        local_tmr_voter(982)  <=    (tmr_registers(0)(982) and tmr_registers(1)(982)) or                                                             
                            (tmr_registers(1)(982) and tmr_registers(2)(982)) or                                                             
                            (tmr_registers(0)(982) and tmr_registers(2)(982));                                                               
                                                                                                                                         
        local_tmr_voter(983)  <=    (tmr_registers(0)(983) and tmr_registers(1)(983)) or                                                             
                            (tmr_registers(1)(983) and tmr_registers(2)(983)) or                                                             
                            (tmr_registers(0)(983) and tmr_registers(2)(983));                                                               
                                                                                                                                         
        local_tmr_voter(984)  <=    (tmr_registers(0)(984) and tmr_registers(1)(984)) or                                                             
                            (tmr_registers(1)(984) and tmr_registers(2)(984)) or                                                             
                            (tmr_registers(0)(984) and tmr_registers(2)(984));                                                               
                                                                                                                                         
        local_tmr_voter(985)  <=    (tmr_registers(0)(985) and tmr_registers(1)(985)) or                                                             
                            (tmr_registers(1)(985) and tmr_registers(2)(985)) or                                                             
                            (tmr_registers(0)(985) and tmr_registers(2)(985));                                                               
                                                                                                                                         
        local_tmr_voter(986)  <=    (tmr_registers(0)(986) and tmr_registers(1)(986)) or                                                             
                            (tmr_registers(1)(986) and tmr_registers(2)(986)) or                                                             
                            (tmr_registers(0)(986) and tmr_registers(2)(986));                                                               
                                                                                                                                         
        local_tmr_voter(987)  <=    (tmr_registers(0)(987) and tmr_registers(1)(987)) or                                                             
                            (tmr_registers(1)(987) and tmr_registers(2)(987)) or                                                             
                            (tmr_registers(0)(987) and tmr_registers(2)(987));                                                               
                                                                                                                                         
        local_tmr_voter(988)  <=    (tmr_registers(0)(988) and tmr_registers(1)(988)) or                                                             
                            (tmr_registers(1)(988) and tmr_registers(2)(988)) or                                                             
                            (tmr_registers(0)(988) and tmr_registers(2)(988));                                                               
                                                                                                                                         
        local_tmr_voter(989)  <=    (tmr_registers(0)(989) and tmr_registers(1)(989)) or                                                             
                            (tmr_registers(1)(989) and tmr_registers(2)(989)) or                                                             
                            (tmr_registers(0)(989) and tmr_registers(2)(989));                                                               
                                                                                                                                         
        local_tmr_voter(990)  <=    (tmr_registers(0)(990) and tmr_registers(1)(990)) or                                                             
                            (tmr_registers(1)(990) and tmr_registers(2)(990)) or                                                             
                            (tmr_registers(0)(990) and tmr_registers(2)(990));                                                               
                                                                                                                                         
        local_tmr_voter(991)  <=    (tmr_registers(0)(991) and tmr_registers(1)(991)) or                                                             
                            (tmr_registers(1)(991) and tmr_registers(2)(991)) or                                                             
                            (tmr_registers(0)(991) and tmr_registers(2)(991));                                                               
                                                                                                                                         
        local_tmr_voter(992)  <=    (tmr_registers(0)(992) and tmr_registers(1)(992)) or                                                             
                            (tmr_registers(1)(992) and tmr_registers(2)(992)) or                                                             
                            (tmr_registers(0)(992) and tmr_registers(2)(992));                                                               
                                                                                                                                         
        local_tmr_voter(993)  <=    (tmr_registers(0)(993) and tmr_registers(1)(993)) or                                                             
                            (tmr_registers(1)(993) and tmr_registers(2)(993)) or                                                             
                            (tmr_registers(0)(993) and tmr_registers(2)(993));                                                               
                                                                                                                                         
        local_tmr_voter(994)  <=    (tmr_registers(0)(994) and tmr_registers(1)(994)) or                                                             
                            (tmr_registers(1)(994) and tmr_registers(2)(994)) or                                                             
                            (tmr_registers(0)(994) and tmr_registers(2)(994));                                                               
                                                                                                                                         
        local_tmr_voter(995)  <=    (tmr_registers(0)(995) and tmr_registers(1)(995)) or                                                             
                            (tmr_registers(1)(995) and tmr_registers(2)(995)) or                                                             
                            (tmr_registers(0)(995) and tmr_registers(2)(995));                                                               
                                                                                                                                         
        local_tmr_voter(996)  <=    (tmr_registers(0)(996) and tmr_registers(1)(996)) or                                                             
                            (tmr_registers(1)(996) and tmr_registers(2)(996)) or                                                             
                            (tmr_registers(0)(996) and tmr_registers(2)(996));                                                               
                                                                                                                                         
        local_tmr_voter(997)  <=    (tmr_registers(0)(997) and tmr_registers(1)(997)) or                                                             
                            (tmr_registers(1)(997) and tmr_registers(2)(997)) or                                                             
                            (tmr_registers(0)(997) and tmr_registers(2)(997));                                                               
                                                                                                                                         
        local_tmr_voter(998)  <=    (tmr_registers(0)(998) and tmr_registers(1)(998)) or                                                             
                            (tmr_registers(1)(998) and tmr_registers(2)(998)) or                                                             
                            (tmr_registers(0)(998) and tmr_registers(2)(998));                                                               
                                                                                                                                         
        local_tmr_voter(999)  <=    (tmr_registers(0)(999) and tmr_registers(1)(999)) or                                                             
                            (tmr_registers(1)(999) and tmr_registers(2)(999)) or                                                             
                            (tmr_registers(0)(999) and tmr_registers(2)(999));                                                               
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Outputs                                                                                                                           
    ------------------------------------------                                                                                           
                                                                                                                                         
    data_out(0) <= local_tmr_voter(nb_reg-4);                                                                                                  
    data_out(1) <= local_tmr_voter(nb_reg-3);                                                                                                  
    data_out(2) <= local_tmr_voter(nb_reg-2);                                                                                                  
    data_out(3) <= local_tmr_voter(nb_reg-1);                                                                                                  
                                                                                                                                         
                                                                                                                                         
end generate LOCAL_TMR_MITIGATION;                                                                                                       
                                                                                                                                         
----------------------------------------------------------------------------------------------------------------------------             
--                                                                                                                                       
--                                                                                                                                       
--              Global TMR                                                                                                               
--                                                                                                                                       
--                                                                                                                                       
----------------------------------------------------------------------------------------------------------------------------             
                                                                                                                                         
GLOBAL_TMR_MITIGATION: if USE_MITIGATION=2 generate                                                                                      
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Input                                                                                                                             
    ------------------------------------------                                                                                           
                                                                                                                                         
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Combinatiorial + Registers                                                                                                        
    ------------------------------------------                                                                                           
    process(clk)                                                                                                                         
    begin                                                                                                                                
                                                                                                                                         
        if rising_edge(clk) then                                                                                                         
                                                                                                                                         
                tmr_registers(0)(1)    <= not(global_tmr_voter(0)(0));                                                             
                tmr_registers(1)(1)    <= not(global_tmr_voter(1)(0));                                                             
                tmr_registers(2)(1)    <= not(global_tmr_voter(2)(0));                                                             
 
                tmr_registers(0)(2)    <= not(global_tmr_voter(0)(1));                                                             
                tmr_registers(1)(2)    <= not(global_tmr_voter(1)(1));                                                             
                tmr_registers(2)(2)    <= not(global_tmr_voter(2)(1));                                                             
 
                tmr_registers(0)(3)    <= not(global_tmr_voter(0)(2));                                                             
                tmr_registers(1)(3)    <= not(global_tmr_voter(1)(2));                                                             
                tmr_registers(2)(3)    <= not(global_tmr_voter(2)(2));                                                             
 
                tmr_registers(0)(4)    <= not(global_tmr_voter(0)(3));                                                             
                tmr_registers(1)(4)    <= not(global_tmr_voter(1)(3));                                                             
                tmr_registers(2)(4)    <= not(global_tmr_voter(2)(3));                                                             
 
                tmr_registers(0)(5)    <= not(global_tmr_voter(0)(4));                                                             
                tmr_registers(1)(5)    <= not(global_tmr_voter(1)(4));                                                             
                tmr_registers(2)(5)    <= not(global_tmr_voter(2)(4));                                                             
 
                tmr_registers(0)(6)    <= not(global_tmr_voter(0)(5));                                                             
                tmr_registers(1)(6)    <= not(global_tmr_voter(1)(5));                                                             
                tmr_registers(2)(6)    <= not(global_tmr_voter(2)(5));                                                             
 
                tmr_registers(0)(7)    <= not(global_tmr_voter(0)(6));                                                             
                tmr_registers(1)(7)    <= not(global_tmr_voter(1)(6));                                                             
                tmr_registers(2)(7)    <= not(global_tmr_voter(2)(6));                                                             
 
                tmr_registers(0)(8)    <= not(global_tmr_voter(0)(7));                                                             
                tmr_registers(1)(8)    <= not(global_tmr_voter(1)(7));                                                             
                tmr_registers(2)(8)    <= not(global_tmr_voter(2)(7));                                                             
 
                tmr_registers(0)(9)    <= not(global_tmr_voter(0)(8));                                                             
                tmr_registers(1)(9)    <= not(global_tmr_voter(1)(8));                                                             
                tmr_registers(2)(9)    <= not(global_tmr_voter(2)(8));                                                             
 
                tmr_registers(0)(10)    <= not(global_tmr_voter(0)(9));                                                             
                tmr_registers(1)(10)    <= not(global_tmr_voter(1)(9));                                                             
                tmr_registers(2)(10)    <= not(global_tmr_voter(2)(9));                                                             
 
                tmr_registers(0)(11)    <= not(global_tmr_voter(0)(10));                                                             
                tmr_registers(1)(11)    <= not(global_tmr_voter(1)(10));                                                             
                tmr_registers(2)(11)    <= not(global_tmr_voter(2)(10));                                                             
 
                tmr_registers(0)(12)    <= not(global_tmr_voter(0)(11));                                                             
                tmr_registers(1)(12)    <= not(global_tmr_voter(1)(11));                                                             
                tmr_registers(2)(12)    <= not(global_tmr_voter(2)(11));                                                             
 
                tmr_registers(0)(13)    <= not(global_tmr_voter(0)(12));                                                             
                tmr_registers(1)(13)    <= not(global_tmr_voter(1)(12));                                                             
                tmr_registers(2)(13)    <= not(global_tmr_voter(2)(12));                                                             
 
                tmr_registers(0)(14)    <= not(global_tmr_voter(0)(13));                                                             
                tmr_registers(1)(14)    <= not(global_tmr_voter(1)(13));                                                             
                tmr_registers(2)(14)    <= not(global_tmr_voter(2)(13));                                                             
 
                tmr_registers(0)(15)    <= not(global_tmr_voter(0)(14));                                                             
                tmr_registers(1)(15)    <= not(global_tmr_voter(1)(14));                                                             
                tmr_registers(2)(15)    <= not(global_tmr_voter(2)(14));                                                             
 
                tmr_registers(0)(16)    <= not(global_tmr_voter(0)(15));                                                             
                tmr_registers(1)(16)    <= not(global_tmr_voter(1)(15));                                                             
                tmr_registers(2)(16)    <= not(global_tmr_voter(2)(15));                                                             
 
                tmr_registers(0)(17)    <= not(global_tmr_voter(0)(16));                                                             
                tmr_registers(1)(17)    <= not(global_tmr_voter(1)(16));                                                             
                tmr_registers(2)(17)    <= not(global_tmr_voter(2)(16));                                                             
 
                tmr_registers(0)(18)    <= not(global_tmr_voter(0)(17));                                                             
                tmr_registers(1)(18)    <= not(global_tmr_voter(1)(17));                                                             
                tmr_registers(2)(18)    <= not(global_tmr_voter(2)(17));                                                             
 
                tmr_registers(0)(19)    <= not(global_tmr_voter(0)(18));                                                             
                tmr_registers(1)(19)    <= not(global_tmr_voter(1)(18));                                                             
                tmr_registers(2)(19)    <= not(global_tmr_voter(2)(18));                                                             
 
                tmr_registers(0)(20)    <= not(global_tmr_voter(0)(19));                                                             
                tmr_registers(1)(20)    <= not(global_tmr_voter(1)(19));                                                             
                tmr_registers(2)(20)    <= not(global_tmr_voter(2)(19));                                                             
 
                tmr_registers(0)(21)    <= not(global_tmr_voter(0)(20));                                                             
                tmr_registers(1)(21)    <= not(global_tmr_voter(1)(20));                                                             
                tmr_registers(2)(21)    <= not(global_tmr_voter(2)(20));                                                             
 
                tmr_registers(0)(22)    <= not(global_tmr_voter(0)(21));                                                             
                tmr_registers(1)(22)    <= not(global_tmr_voter(1)(21));                                                             
                tmr_registers(2)(22)    <= not(global_tmr_voter(2)(21));                                                             
 
                tmr_registers(0)(23)    <= not(global_tmr_voter(0)(22));                                                             
                tmr_registers(1)(23)    <= not(global_tmr_voter(1)(22));                                                             
                tmr_registers(2)(23)    <= not(global_tmr_voter(2)(22));                                                             
 
                tmr_registers(0)(24)    <= not(global_tmr_voter(0)(23));                                                             
                tmr_registers(1)(24)    <= not(global_tmr_voter(1)(23));                                                             
                tmr_registers(2)(24)    <= not(global_tmr_voter(2)(23));                                                             
 
                tmr_registers(0)(25)    <= not(global_tmr_voter(0)(24));                                                             
                tmr_registers(1)(25)    <= not(global_tmr_voter(1)(24));                                                             
                tmr_registers(2)(25)    <= not(global_tmr_voter(2)(24));                                                             
 
                tmr_registers(0)(26)    <= not(global_tmr_voter(0)(25));                                                             
                tmr_registers(1)(26)    <= not(global_tmr_voter(1)(25));                                                             
                tmr_registers(2)(26)    <= not(global_tmr_voter(2)(25));                                                             
 
                tmr_registers(0)(27)    <= not(global_tmr_voter(0)(26));                                                             
                tmr_registers(1)(27)    <= not(global_tmr_voter(1)(26));                                                             
                tmr_registers(2)(27)    <= not(global_tmr_voter(2)(26));                                                             
 
                tmr_registers(0)(28)    <= not(global_tmr_voter(0)(27));                                                             
                tmr_registers(1)(28)    <= not(global_tmr_voter(1)(27));                                                             
                tmr_registers(2)(28)    <= not(global_tmr_voter(2)(27));                                                             
 
                tmr_registers(0)(29)    <= not(global_tmr_voter(0)(28));                                                             
                tmr_registers(1)(29)    <= not(global_tmr_voter(1)(28));                                                             
                tmr_registers(2)(29)    <= not(global_tmr_voter(2)(28));                                                             
 
                tmr_registers(0)(30)    <= not(global_tmr_voter(0)(29));                                                             
                tmr_registers(1)(30)    <= not(global_tmr_voter(1)(29));                                                             
                tmr_registers(2)(30)    <= not(global_tmr_voter(2)(29));                                                             
 
                tmr_registers(0)(31)    <= not(global_tmr_voter(0)(30));                                                             
                tmr_registers(1)(31)    <= not(global_tmr_voter(1)(30));                                                             
                tmr_registers(2)(31)    <= not(global_tmr_voter(2)(30));                                                             
 
                tmr_registers(0)(32)    <= not(global_tmr_voter(0)(31));                                                             
                tmr_registers(1)(32)    <= not(global_tmr_voter(1)(31));                                                             
                tmr_registers(2)(32)    <= not(global_tmr_voter(2)(31));                                                             
 
                tmr_registers(0)(33)    <= not(global_tmr_voter(0)(32));                                                             
                tmr_registers(1)(33)    <= not(global_tmr_voter(1)(32));                                                             
                tmr_registers(2)(33)    <= not(global_tmr_voter(2)(32));                                                             
 
                tmr_registers(0)(34)    <= not(global_tmr_voter(0)(33));                                                             
                tmr_registers(1)(34)    <= not(global_tmr_voter(1)(33));                                                             
                tmr_registers(2)(34)    <= not(global_tmr_voter(2)(33));                                                             
 
                tmr_registers(0)(35)    <= not(global_tmr_voter(0)(34));                                                             
                tmr_registers(1)(35)    <= not(global_tmr_voter(1)(34));                                                             
                tmr_registers(2)(35)    <= not(global_tmr_voter(2)(34));                                                             
 
                tmr_registers(0)(36)    <= not(global_tmr_voter(0)(35));                                                             
                tmr_registers(1)(36)    <= not(global_tmr_voter(1)(35));                                                             
                tmr_registers(2)(36)    <= not(global_tmr_voter(2)(35));                                                             
 
                tmr_registers(0)(37)    <= not(global_tmr_voter(0)(36));                                                             
                tmr_registers(1)(37)    <= not(global_tmr_voter(1)(36));                                                             
                tmr_registers(2)(37)    <= not(global_tmr_voter(2)(36));                                                             
 
                tmr_registers(0)(38)    <= not(global_tmr_voter(0)(37));                                                             
                tmr_registers(1)(38)    <= not(global_tmr_voter(1)(37));                                                             
                tmr_registers(2)(38)    <= not(global_tmr_voter(2)(37));                                                             
 
                tmr_registers(0)(39)    <= not(global_tmr_voter(0)(38));                                                             
                tmr_registers(1)(39)    <= not(global_tmr_voter(1)(38));                                                             
                tmr_registers(2)(39)    <= not(global_tmr_voter(2)(38));                                                             
 
                tmr_registers(0)(40)    <= not(global_tmr_voter(0)(39));                                                             
                tmr_registers(1)(40)    <= not(global_tmr_voter(1)(39));                                                             
                tmr_registers(2)(40)    <= not(global_tmr_voter(2)(39));                                                             
 
                tmr_registers(0)(41)    <= not(global_tmr_voter(0)(40));                                                             
                tmr_registers(1)(41)    <= not(global_tmr_voter(1)(40));                                                             
                tmr_registers(2)(41)    <= not(global_tmr_voter(2)(40));                                                             
 
                tmr_registers(0)(42)    <= not(global_tmr_voter(0)(41));                                                             
                tmr_registers(1)(42)    <= not(global_tmr_voter(1)(41));                                                             
                tmr_registers(2)(42)    <= not(global_tmr_voter(2)(41));                                                             
 
                tmr_registers(0)(43)    <= not(global_tmr_voter(0)(42));                                                             
                tmr_registers(1)(43)    <= not(global_tmr_voter(1)(42));                                                             
                tmr_registers(2)(43)    <= not(global_tmr_voter(2)(42));                                                             
 
                tmr_registers(0)(44)    <= not(global_tmr_voter(0)(43));                                                             
                tmr_registers(1)(44)    <= not(global_tmr_voter(1)(43));                                                             
                tmr_registers(2)(44)    <= not(global_tmr_voter(2)(43));                                                             
 
                tmr_registers(0)(45)    <= not(global_tmr_voter(0)(44));                                                             
                tmr_registers(1)(45)    <= not(global_tmr_voter(1)(44));                                                             
                tmr_registers(2)(45)    <= not(global_tmr_voter(2)(44));                                                             
 
                tmr_registers(0)(46)    <= not(global_tmr_voter(0)(45));                                                             
                tmr_registers(1)(46)    <= not(global_tmr_voter(1)(45));                                                             
                tmr_registers(2)(46)    <= not(global_tmr_voter(2)(45));                                                             
 
                tmr_registers(0)(47)    <= not(global_tmr_voter(0)(46));                                                             
                tmr_registers(1)(47)    <= not(global_tmr_voter(1)(46));                                                             
                tmr_registers(2)(47)    <= not(global_tmr_voter(2)(46));                                                             
 
                tmr_registers(0)(48)    <= not(global_tmr_voter(0)(47));                                                             
                tmr_registers(1)(48)    <= not(global_tmr_voter(1)(47));                                                             
                tmr_registers(2)(48)    <= not(global_tmr_voter(2)(47));                                                             
 
                tmr_registers(0)(49)    <= not(global_tmr_voter(0)(48));                                                             
                tmr_registers(1)(49)    <= not(global_tmr_voter(1)(48));                                                             
                tmr_registers(2)(49)    <= not(global_tmr_voter(2)(48));                                                             
 
                tmr_registers(0)(50)    <= not(global_tmr_voter(0)(49));                                                             
                tmr_registers(1)(50)    <= not(global_tmr_voter(1)(49));                                                             
                tmr_registers(2)(50)    <= not(global_tmr_voter(2)(49));                                                             
 
                tmr_registers(0)(51)    <= not(global_tmr_voter(0)(50));                                                             
                tmr_registers(1)(51)    <= not(global_tmr_voter(1)(50));                                                             
                tmr_registers(2)(51)    <= not(global_tmr_voter(2)(50));                                                             
 
                tmr_registers(0)(52)    <= not(global_tmr_voter(0)(51));                                                             
                tmr_registers(1)(52)    <= not(global_tmr_voter(1)(51));                                                             
                tmr_registers(2)(52)    <= not(global_tmr_voter(2)(51));                                                             
 
                tmr_registers(0)(53)    <= not(global_tmr_voter(0)(52));                                                             
                tmr_registers(1)(53)    <= not(global_tmr_voter(1)(52));                                                             
                tmr_registers(2)(53)    <= not(global_tmr_voter(2)(52));                                                             
 
                tmr_registers(0)(54)    <= not(global_tmr_voter(0)(53));                                                             
                tmr_registers(1)(54)    <= not(global_tmr_voter(1)(53));                                                             
                tmr_registers(2)(54)    <= not(global_tmr_voter(2)(53));                                                             
 
                tmr_registers(0)(55)    <= not(global_tmr_voter(0)(54));                                                             
                tmr_registers(1)(55)    <= not(global_tmr_voter(1)(54));                                                             
                tmr_registers(2)(55)    <= not(global_tmr_voter(2)(54));                                                             
 
                tmr_registers(0)(56)    <= not(global_tmr_voter(0)(55));                                                             
                tmr_registers(1)(56)    <= not(global_tmr_voter(1)(55));                                                             
                tmr_registers(2)(56)    <= not(global_tmr_voter(2)(55));                                                             
 
                tmr_registers(0)(57)    <= not(global_tmr_voter(0)(56));                                                             
                tmr_registers(1)(57)    <= not(global_tmr_voter(1)(56));                                                             
                tmr_registers(2)(57)    <= not(global_tmr_voter(2)(56));                                                             
 
                tmr_registers(0)(58)    <= not(global_tmr_voter(0)(57));                                                             
                tmr_registers(1)(58)    <= not(global_tmr_voter(1)(57));                                                             
                tmr_registers(2)(58)    <= not(global_tmr_voter(2)(57));                                                             
 
                tmr_registers(0)(59)    <= not(global_tmr_voter(0)(58));                                                             
                tmr_registers(1)(59)    <= not(global_tmr_voter(1)(58));                                                             
                tmr_registers(2)(59)    <= not(global_tmr_voter(2)(58));                                                             
 
                tmr_registers(0)(60)    <= not(global_tmr_voter(0)(59));                                                             
                tmr_registers(1)(60)    <= not(global_tmr_voter(1)(59));                                                             
                tmr_registers(2)(60)    <= not(global_tmr_voter(2)(59));                                                             
 
                tmr_registers(0)(61)    <= not(global_tmr_voter(0)(60));                                                             
                tmr_registers(1)(61)    <= not(global_tmr_voter(1)(60));                                                             
                tmr_registers(2)(61)    <= not(global_tmr_voter(2)(60));                                                             
 
                tmr_registers(0)(62)    <= not(global_tmr_voter(0)(61));                                                             
                tmr_registers(1)(62)    <= not(global_tmr_voter(1)(61));                                                             
                tmr_registers(2)(62)    <= not(global_tmr_voter(2)(61));                                                             
 
                tmr_registers(0)(63)    <= not(global_tmr_voter(0)(62));                                                             
                tmr_registers(1)(63)    <= not(global_tmr_voter(1)(62));                                                             
                tmr_registers(2)(63)    <= not(global_tmr_voter(2)(62));                                                             
 
                tmr_registers(0)(64)    <= not(global_tmr_voter(0)(63));                                                             
                tmr_registers(1)(64)    <= not(global_tmr_voter(1)(63));                                                             
                tmr_registers(2)(64)    <= not(global_tmr_voter(2)(63));                                                             
 
                tmr_registers(0)(65)    <= not(global_tmr_voter(0)(64));                                                             
                tmr_registers(1)(65)    <= not(global_tmr_voter(1)(64));                                                             
                tmr_registers(2)(65)    <= not(global_tmr_voter(2)(64));                                                             
 
                tmr_registers(0)(66)    <= not(global_tmr_voter(0)(65));                                                             
                tmr_registers(1)(66)    <= not(global_tmr_voter(1)(65));                                                             
                tmr_registers(2)(66)    <= not(global_tmr_voter(2)(65));                                                             
 
                tmr_registers(0)(67)    <= not(global_tmr_voter(0)(66));                                                             
                tmr_registers(1)(67)    <= not(global_tmr_voter(1)(66));                                                             
                tmr_registers(2)(67)    <= not(global_tmr_voter(2)(66));                                                             
 
                tmr_registers(0)(68)    <= not(global_tmr_voter(0)(67));                                                             
                tmr_registers(1)(68)    <= not(global_tmr_voter(1)(67));                                                             
                tmr_registers(2)(68)    <= not(global_tmr_voter(2)(67));                                                             
 
                tmr_registers(0)(69)    <= not(global_tmr_voter(0)(68));                                                             
                tmr_registers(1)(69)    <= not(global_tmr_voter(1)(68));                                                             
                tmr_registers(2)(69)    <= not(global_tmr_voter(2)(68));                                                             
 
                tmr_registers(0)(70)    <= not(global_tmr_voter(0)(69));                                                             
                tmr_registers(1)(70)    <= not(global_tmr_voter(1)(69));                                                             
                tmr_registers(2)(70)    <= not(global_tmr_voter(2)(69));                                                             
 
                tmr_registers(0)(71)    <= not(global_tmr_voter(0)(70));                                                             
                tmr_registers(1)(71)    <= not(global_tmr_voter(1)(70));                                                             
                tmr_registers(2)(71)    <= not(global_tmr_voter(2)(70));                                                             
 
                tmr_registers(0)(72)    <= not(global_tmr_voter(0)(71));                                                             
                tmr_registers(1)(72)    <= not(global_tmr_voter(1)(71));                                                             
                tmr_registers(2)(72)    <= not(global_tmr_voter(2)(71));                                                             
 
                tmr_registers(0)(73)    <= not(global_tmr_voter(0)(72));                                                             
                tmr_registers(1)(73)    <= not(global_tmr_voter(1)(72));                                                             
                tmr_registers(2)(73)    <= not(global_tmr_voter(2)(72));                                                             
 
                tmr_registers(0)(74)    <= not(global_tmr_voter(0)(73));                                                             
                tmr_registers(1)(74)    <= not(global_tmr_voter(1)(73));                                                             
                tmr_registers(2)(74)    <= not(global_tmr_voter(2)(73));                                                             
 
                tmr_registers(0)(75)    <= not(global_tmr_voter(0)(74));                                                             
                tmr_registers(1)(75)    <= not(global_tmr_voter(1)(74));                                                             
                tmr_registers(2)(75)    <= not(global_tmr_voter(2)(74));                                                             
 
                tmr_registers(0)(76)    <= not(global_tmr_voter(0)(75));                                                             
                tmr_registers(1)(76)    <= not(global_tmr_voter(1)(75));                                                             
                tmr_registers(2)(76)    <= not(global_tmr_voter(2)(75));                                                             
 
                tmr_registers(0)(77)    <= not(global_tmr_voter(0)(76));                                                             
                tmr_registers(1)(77)    <= not(global_tmr_voter(1)(76));                                                             
                tmr_registers(2)(77)    <= not(global_tmr_voter(2)(76));                                                             
 
                tmr_registers(0)(78)    <= not(global_tmr_voter(0)(77));                                                             
                tmr_registers(1)(78)    <= not(global_tmr_voter(1)(77));                                                             
                tmr_registers(2)(78)    <= not(global_tmr_voter(2)(77));                                                             
 
                tmr_registers(0)(79)    <= not(global_tmr_voter(0)(78));                                                             
                tmr_registers(1)(79)    <= not(global_tmr_voter(1)(78));                                                             
                tmr_registers(2)(79)    <= not(global_tmr_voter(2)(78));                                                             
 
                tmr_registers(0)(80)    <= not(global_tmr_voter(0)(79));                                                             
                tmr_registers(1)(80)    <= not(global_tmr_voter(1)(79));                                                             
                tmr_registers(2)(80)    <= not(global_tmr_voter(2)(79));                                                             
 
                tmr_registers(0)(81)    <= not(global_tmr_voter(0)(80));                                                             
                tmr_registers(1)(81)    <= not(global_tmr_voter(1)(80));                                                             
                tmr_registers(2)(81)    <= not(global_tmr_voter(2)(80));                                                             
 
                tmr_registers(0)(82)    <= not(global_tmr_voter(0)(81));                                                             
                tmr_registers(1)(82)    <= not(global_tmr_voter(1)(81));                                                             
                tmr_registers(2)(82)    <= not(global_tmr_voter(2)(81));                                                             
 
                tmr_registers(0)(83)    <= not(global_tmr_voter(0)(82));                                                             
                tmr_registers(1)(83)    <= not(global_tmr_voter(1)(82));                                                             
                tmr_registers(2)(83)    <= not(global_tmr_voter(2)(82));                                                             
 
                tmr_registers(0)(84)    <= not(global_tmr_voter(0)(83));                                                             
                tmr_registers(1)(84)    <= not(global_tmr_voter(1)(83));                                                             
                tmr_registers(2)(84)    <= not(global_tmr_voter(2)(83));                                                             
 
                tmr_registers(0)(85)    <= not(global_tmr_voter(0)(84));                                                             
                tmr_registers(1)(85)    <= not(global_tmr_voter(1)(84));                                                             
                tmr_registers(2)(85)    <= not(global_tmr_voter(2)(84));                                                             
 
                tmr_registers(0)(86)    <= not(global_tmr_voter(0)(85));                                                             
                tmr_registers(1)(86)    <= not(global_tmr_voter(1)(85));                                                             
                tmr_registers(2)(86)    <= not(global_tmr_voter(2)(85));                                                             
 
                tmr_registers(0)(87)    <= not(global_tmr_voter(0)(86));                                                             
                tmr_registers(1)(87)    <= not(global_tmr_voter(1)(86));                                                             
                tmr_registers(2)(87)    <= not(global_tmr_voter(2)(86));                                                             
 
                tmr_registers(0)(88)    <= not(global_tmr_voter(0)(87));                                                             
                tmr_registers(1)(88)    <= not(global_tmr_voter(1)(87));                                                             
                tmr_registers(2)(88)    <= not(global_tmr_voter(2)(87));                                                             
 
                tmr_registers(0)(89)    <= not(global_tmr_voter(0)(88));                                                             
                tmr_registers(1)(89)    <= not(global_tmr_voter(1)(88));                                                             
                tmr_registers(2)(89)    <= not(global_tmr_voter(2)(88));                                                             
 
                tmr_registers(0)(90)    <= not(global_tmr_voter(0)(89));                                                             
                tmr_registers(1)(90)    <= not(global_tmr_voter(1)(89));                                                             
                tmr_registers(2)(90)    <= not(global_tmr_voter(2)(89));                                                             
 
                tmr_registers(0)(91)    <= not(global_tmr_voter(0)(90));                                                             
                tmr_registers(1)(91)    <= not(global_tmr_voter(1)(90));                                                             
                tmr_registers(2)(91)    <= not(global_tmr_voter(2)(90));                                                             
 
                tmr_registers(0)(92)    <= not(global_tmr_voter(0)(91));                                                             
                tmr_registers(1)(92)    <= not(global_tmr_voter(1)(91));                                                             
                tmr_registers(2)(92)    <= not(global_tmr_voter(2)(91));                                                             
 
                tmr_registers(0)(93)    <= not(global_tmr_voter(0)(92));                                                             
                tmr_registers(1)(93)    <= not(global_tmr_voter(1)(92));                                                             
                tmr_registers(2)(93)    <= not(global_tmr_voter(2)(92));                                                             
 
                tmr_registers(0)(94)    <= not(global_tmr_voter(0)(93));                                                             
                tmr_registers(1)(94)    <= not(global_tmr_voter(1)(93));                                                             
                tmr_registers(2)(94)    <= not(global_tmr_voter(2)(93));                                                             
 
                tmr_registers(0)(95)    <= not(global_tmr_voter(0)(94));                                                             
                tmr_registers(1)(95)    <= not(global_tmr_voter(1)(94));                                                             
                tmr_registers(2)(95)    <= not(global_tmr_voter(2)(94));                                                             
 
                tmr_registers(0)(96)    <= not(global_tmr_voter(0)(95));                                                             
                tmr_registers(1)(96)    <= not(global_tmr_voter(1)(95));                                                             
                tmr_registers(2)(96)    <= not(global_tmr_voter(2)(95));                                                             
 
                tmr_registers(0)(97)    <= not(global_tmr_voter(0)(96));                                                             
                tmr_registers(1)(97)    <= not(global_tmr_voter(1)(96));                                                             
                tmr_registers(2)(97)    <= not(global_tmr_voter(2)(96));                                                             
 
                tmr_registers(0)(98)    <= not(global_tmr_voter(0)(97));                                                             
                tmr_registers(1)(98)    <= not(global_tmr_voter(1)(97));                                                             
                tmr_registers(2)(98)    <= not(global_tmr_voter(2)(97));                                                             
 
                tmr_registers(0)(99)    <= not(global_tmr_voter(0)(98));                                                             
                tmr_registers(1)(99)    <= not(global_tmr_voter(1)(98));                                                             
                tmr_registers(2)(99)    <= not(global_tmr_voter(2)(98));                                                             
 
                tmr_registers(0)(100)    <= not(global_tmr_voter(0)(99));                                                             
                tmr_registers(1)(100)    <= not(global_tmr_voter(1)(99));                                                             
                tmr_registers(2)(100)    <= not(global_tmr_voter(2)(99));                                                             
 
                tmr_registers(0)(101)    <= not(global_tmr_voter(0)(100));                                                             
                tmr_registers(1)(101)    <= not(global_tmr_voter(1)(100));                                                             
                tmr_registers(2)(101)    <= not(global_tmr_voter(2)(100));                                                             
 
                tmr_registers(0)(102)    <= not(global_tmr_voter(0)(101));                                                             
                tmr_registers(1)(102)    <= not(global_tmr_voter(1)(101));                                                             
                tmr_registers(2)(102)    <= not(global_tmr_voter(2)(101));                                                             
 
                tmr_registers(0)(103)    <= not(global_tmr_voter(0)(102));                                                             
                tmr_registers(1)(103)    <= not(global_tmr_voter(1)(102));                                                             
                tmr_registers(2)(103)    <= not(global_tmr_voter(2)(102));                                                             
 
                tmr_registers(0)(104)    <= not(global_tmr_voter(0)(103));                                                             
                tmr_registers(1)(104)    <= not(global_tmr_voter(1)(103));                                                             
                tmr_registers(2)(104)    <= not(global_tmr_voter(2)(103));                                                             
 
                tmr_registers(0)(105)    <= not(global_tmr_voter(0)(104));                                                             
                tmr_registers(1)(105)    <= not(global_tmr_voter(1)(104));                                                             
                tmr_registers(2)(105)    <= not(global_tmr_voter(2)(104));                                                             
 
                tmr_registers(0)(106)    <= not(global_tmr_voter(0)(105));                                                             
                tmr_registers(1)(106)    <= not(global_tmr_voter(1)(105));                                                             
                tmr_registers(2)(106)    <= not(global_tmr_voter(2)(105));                                                             
 
                tmr_registers(0)(107)    <= not(global_tmr_voter(0)(106));                                                             
                tmr_registers(1)(107)    <= not(global_tmr_voter(1)(106));                                                             
                tmr_registers(2)(107)    <= not(global_tmr_voter(2)(106));                                                             
 
                tmr_registers(0)(108)    <= not(global_tmr_voter(0)(107));                                                             
                tmr_registers(1)(108)    <= not(global_tmr_voter(1)(107));                                                             
                tmr_registers(2)(108)    <= not(global_tmr_voter(2)(107));                                                             
 
                tmr_registers(0)(109)    <= not(global_tmr_voter(0)(108));                                                             
                tmr_registers(1)(109)    <= not(global_tmr_voter(1)(108));                                                             
                tmr_registers(2)(109)    <= not(global_tmr_voter(2)(108));                                                             
 
                tmr_registers(0)(110)    <= not(global_tmr_voter(0)(109));                                                             
                tmr_registers(1)(110)    <= not(global_tmr_voter(1)(109));                                                             
                tmr_registers(2)(110)    <= not(global_tmr_voter(2)(109));                                                             
 
                tmr_registers(0)(111)    <= not(global_tmr_voter(0)(110));                                                             
                tmr_registers(1)(111)    <= not(global_tmr_voter(1)(110));                                                             
                tmr_registers(2)(111)    <= not(global_tmr_voter(2)(110));                                                             
 
                tmr_registers(0)(112)    <= not(global_tmr_voter(0)(111));                                                             
                tmr_registers(1)(112)    <= not(global_tmr_voter(1)(111));                                                             
                tmr_registers(2)(112)    <= not(global_tmr_voter(2)(111));                                                             
 
                tmr_registers(0)(113)    <= not(global_tmr_voter(0)(112));                                                             
                tmr_registers(1)(113)    <= not(global_tmr_voter(1)(112));                                                             
                tmr_registers(2)(113)    <= not(global_tmr_voter(2)(112));                                                             
 
                tmr_registers(0)(114)    <= not(global_tmr_voter(0)(113));                                                             
                tmr_registers(1)(114)    <= not(global_tmr_voter(1)(113));                                                             
                tmr_registers(2)(114)    <= not(global_tmr_voter(2)(113));                                                             
 
                tmr_registers(0)(115)    <= not(global_tmr_voter(0)(114));                                                             
                tmr_registers(1)(115)    <= not(global_tmr_voter(1)(114));                                                             
                tmr_registers(2)(115)    <= not(global_tmr_voter(2)(114));                                                             
 
                tmr_registers(0)(116)    <= not(global_tmr_voter(0)(115));                                                             
                tmr_registers(1)(116)    <= not(global_tmr_voter(1)(115));                                                             
                tmr_registers(2)(116)    <= not(global_tmr_voter(2)(115));                                                             
 
                tmr_registers(0)(117)    <= not(global_tmr_voter(0)(116));                                                             
                tmr_registers(1)(117)    <= not(global_tmr_voter(1)(116));                                                             
                tmr_registers(2)(117)    <= not(global_tmr_voter(2)(116));                                                             
 
                tmr_registers(0)(118)    <= not(global_tmr_voter(0)(117));                                                             
                tmr_registers(1)(118)    <= not(global_tmr_voter(1)(117));                                                             
                tmr_registers(2)(118)    <= not(global_tmr_voter(2)(117));                                                             
 
                tmr_registers(0)(119)    <= not(global_tmr_voter(0)(118));                                                             
                tmr_registers(1)(119)    <= not(global_tmr_voter(1)(118));                                                             
                tmr_registers(2)(119)    <= not(global_tmr_voter(2)(118));                                                             
 
                tmr_registers(0)(120)    <= not(global_tmr_voter(0)(119));                                                             
                tmr_registers(1)(120)    <= not(global_tmr_voter(1)(119));                                                             
                tmr_registers(2)(120)    <= not(global_tmr_voter(2)(119));                                                             
 
                tmr_registers(0)(121)    <= not(global_tmr_voter(0)(120));                                                             
                tmr_registers(1)(121)    <= not(global_tmr_voter(1)(120));                                                             
                tmr_registers(2)(121)    <= not(global_tmr_voter(2)(120));                                                             
 
                tmr_registers(0)(122)    <= not(global_tmr_voter(0)(121));                                                             
                tmr_registers(1)(122)    <= not(global_tmr_voter(1)(121));                                                             
                tmr_registers(2)(122)    <= not(global_tmr_voter(2)(121));                                                             
 
                tmr_registers(0)(123)    <= not(global_tmr_voter(0)(122));                                                             
                tmr_registers(1)(123)    <= not(global_tmr_voter(1)(122));                                                             
                tmr_registers(2)(123)    <= not(global_tmr_voter(2)(122));                                                             
 
                tmr_registers(0)(124)    <= not(global_tmr_voter(0)(123));                                                             
                tmr_registers(1)(124)    <= not(global_tmr_voter(1)(123));                                                             
                tmr_registers(2)(124)    <= not(global_tmr_voter(2)(123));                                                             
 
                tmr_registers(0)(125)    <= not(global_tmr_voter(0)(124));                                                             
                tmr_registers(1)(125)    <= not(global_tmr_voter(1)(124));                                                             
                tmr_registers(2)(125)    <= not(global_tmr_voter(2)(124));                                                             
 
                tmr_registers(0)(126)    <= not(global_tmr_voter(0)(125));                                                             
                tmr_registers(1)(126)    <= not(global_tmr_voter(1)(125));                                                             
                tmr_registers(2)(126)    <= not(global_tmr_voter(2)(125));                                                             
 
                tmr_registers(0)(127)    <= not(global_tmr_voter(0)(126));                                                             
                tmr_registers(1)(127)    <= not(global_tmr_voter(1)(126));                                                             
                tmr_registers(2)(127)    <= not(global_tmr_voter(2)(126));                                                             
 
                tmr_registers(0)(128)    <= not(global_tmr_voter(0)(127));                                                             
                tmr_registers(1)(128)    <= not(global_tmr_voter(1)(127));                                                             
                tmr_registers(2)(128)    <= not(global_tmr_voter(2)(127));                                                             
 
                tmr_registers(0)(129)    <= not(global_tmr_voter(0)(128));                                                             
                tmr_registers(1)(129)    <= not(global_tmr_voter(1)(128));                                                             
                tmr_registers(2)(129)    <= not(global_tmr_voter(2)(128));                                                             
 
                tmr_registers(0)(130)    <= not(global_tmr_voter(0)(129));                                                             
                tmr_registers(1)(130)    <= not(global_tmr_voter(1)(129));                                                             
                tmr_registers(2)(130)    <= not(global_tmr_voter(2)(129));                                                             
 
                tmr_registers(0)(131)    <= not(global_tmr_voter(0)(130));                                                             
                tmr_registers(1)(131)    <= not(global_tmr_voter(1)(130));                                                             
                tmr_registers(2)(131)    <= not(global_tmr_voter(2)(130));                                                             
 
                tmr_registers(0)(132)    <= not(global_tmr_voter(0)(131));                                                             
                tmr_registers(1)(132)    <= not(global_tmr_voter(1)(131));                                                             
                tmr_registers(2)(132)    <= not(global_tmr_voter(2)(131));                                                             
 
                tmr_registers(0)(133)    <= not(global_tmr_voter(0)(132));                                                             
                tmr_registers(1)(133)    <= not(global_tmr_voter(1)(132));                                                             
                tmr_registers(2)(133)    <= not(global_tmr_voter(2)(132));                                                             
 
                tmr_registers(0)(134)    <= not(global_tmr_voter(0)(133));                                                             
                tmr_registers(1)(134)    <= not(global_tmr_voter(1)(133));                                                             
                tmr_registers(2)(134)    <= not(global_tmr_voter(2)(133));                                                             
 
                tmr_registers(0)(135)    <= not(global_tmr_voter(0)(134));                                                             
                tmr_registers(1)(135)    <= not(global_tmr_voter(1)(134));                                                             
                tmr_registers(2)(135)    <= not(global_tmr_voter(2)(134));                                                             
 
                tmr_registers(0)(136)    <= not(global_tmr_voter(0)(135));                                                             
                tmr_registers(1)(136)    <= not(global_tmr_voter(1)(135));                                                             
                tmr_registers(2)(136)    <= not(global_tmr_voter(2)(135));                                                             
 
                tmr_registers(0)(137)    <= not(global_tmr_voter(0)(136));                                                             
                tmr_registers(1)(137)    <= not(global_tmr_voter(1)(136));                                                             
                tmr_registers(2)(137)    <= not(global_tmr_voter(2)(136));                                                             
 
                tmr_registers(0)(138)    <= not(global_tmr_voter(0)(137));                                                             
                tmr_registers(1)(138)    <= not(global_tmr_voter(1)(137));                                                             
                tmr_registers(2)(138)    <= not(global_tmr_voter(2)(137));                                                             
 
                tmr_registers(0)(139)    <= not(global_tmr_voter(0)(138));                                                             
                tmr_registers(1)(139)    <= not(global_tmr_voter(1)(138));                                                             
                tmr_registers(2)(139)    <= not(global_tmr_voter(2)(138));                                                             
 
                tmr_registers(0)(140)    <= not(global_tmr_voter(0)(139));                                                             
                tmr_registers(1)(140)    <= not(global_tmr_voter(1)(139));                                                             
                tmr_registers(2)(140)    <= not(global_tmr_voter(2)(139));                                                             
 
                tmr_registers(0)(141)    <= not(global_tmr_voter(0)(140));                                                             
                tmr_registers(1)(141)    <= not(global_tmr_voter(1)(140));                                                             
                tmr_registers(2)(141)    <= not(global_tmr_voter(2)(140));                                                             
 
                tmr_registers(0)(142)    <= not(global_tmr_voter(0)(141));                                                             
                tmr_registers(1)(142)    <= not(global_tmr_voter(1)(141));                                                             
                tmr_registers(2)(142)    <= not(global_tmr_voter(2)(141));                                                             
 
                tmr_registers(0)(143)    <= not(global_tmr_voter(0)(142));                                                             
                tmr_registers(1)(143)    <= not(global_tmr_voter(1)(142));                                                             
                tmr_registers(2)(143)    <= not(global_tmr_voter(2)(142));                                                             
 
                tmr_registers(0)(144)    <= not(global_tmr_voter(0)(143));                                                             
                tmr_registers(1)(144)    <= not(global_tmr_voter(1)(143));                                                             
                tmr_registers(2)(144)    <= not(global_tmr_voter(2)(143));                                                             
 
                tmr_registers(0)(145)    <= not(global_tmr_voter(0)(144));                                                             
                tmr_registers(1)(145)    <= not(global_tmr_voter(1)(144));                                                             
                tmr_registers(2)(145)    <= not(global_tmr_voter(2)(144));                                                             
 
                tmr_registers(0)(146)    <= not(global_tmr_voter(0)(145));                                                             
                tmr_registers(1)(146)    <= not(global_tmr_voter(1)(145));                                                             
                tmr_registers(2)(146)    <= not(global_tmr_voter(2)(145));                                                             
 
                tmr_registers(0)(147)    <= not(global_tmr_voter(0)(146));                                                             
                tmr_registers(1)(147)    <= not(global_tmr_voter(1)(146));                                                             
                tmr_registers(2)(147)    <= not(global_tmr_voter(2)(146));                                                             
 
                tmr_registers(0)(148)    <= not(global_tmr_voter(0)(147));                                                             
                tmr_registers(1)(148)    <= not(global_tmr_voter(1)(147));                                                             
                tmr_registers(2)(148)    <= not(global_tmr_voter(2)(147));                                                             
 
                tmr_registers(0)(149)    <= not(global_tmr_voter(0)(148));                                                             
                tmr_registers(1)(149)    <= not(global_tmr_voter(1)(148));                                                             
                tmr_registers(2)(149)    <= not(global_tmr_voter(2)(148));                                                             
 
                tmr_registers(0)(150)    <= not(global_tmr_voter(0)(149));                                                             
                tmr_registers(1)(150)    <= not(global_tmr_voter(1)(149));                                                             
                tmr_registers(2)(150)    <= not(global_tmr_voter(2)(149));                                                             
 
                tmr_registers(0)(151)    <= not(global_tmr_voter(0)(150));                                                             
                tmr_registers(1)(151)    <= not(global_tmr_voter(1)(150));                                                             
                tmr_registers(2)(151)    <= not(global_tmr_voter(2)(150));                                                             
 
                tmr_registers(0)(152)    <= not(global_tmr_voter(0)(151));                                                             
                tmr_registers(1)(152)    <= not(global_tmr_voter(1)(151));                                                             
                tmr_registers(2)(152)    <= not(global_tmr_voter(2)(151));                                                             
 
                tmr_registers(0)(153)    <= not(global_tmr_voter(0)(152));                                                             
                tmr_registers(1)(153)    <= not(global_tmr_voter(1)(152));                                                             
                tmr_registers(2)(153)    <= not(global_tmr_voter(2)(152));                                                             
 
                tmr_registers(0)(154)    <= not(global_tmr_voter(0)(153));                                                             
                tmr_registers(1)(154)    <= not(global_tmr_voter(1)(153));                                                             
                tmr_registers(2)(154)    <= not(global_tmr_voter(2)(153));                                                             
 
                tmr_registers(0)(155)    <= not(global_tmr_voter(0)(154));                                                             
                tmr_registers(1)(155)    <= not(global_tmr_voter(1)(154));                                                             
                tmr_registers(2)(155)    <= not(global_tmr_voter(2)(154));                                                             
 
                tmr_registers(0)(156)    <= not(global_tmr_voter(0)(155));                                                             
                tmr_registers(1)(156)    <= not(global_tmr_voter(1)(155));                                                             
                tmr_registers(2)(156)    <= not(global_tmr_voter(2)(155));                                                             
 
                tmr_registers(0)(157)    <= not(global_tmr_voter(0)(156));                                                             
                tmr_registers(1)(157)    <= not(global_tmr_voter(1)(156));                                                             
                tmr_registers(2)(157)    <= not(global_tmr_voter(2)(156));                                                             
 
                tmr_registers(0)(158)    <= not(global_tmr_voter(0)(157));                                                             
                tmr_registers(1)(158)    <= not(global_tmr_voter(1)(157));                                                             
                tmr_registers(2)(158)    <= not(global_tmr_voter(2)(157));                                                             
 
                tmr_registers(0)(159)    <= not(global_tmr_voter(0)(158));                                                             
                tmr_registers(1)(159)    <= not(global_tmr_voter(1)(158));                                                             
                tmr_registers(2)(159)    <= not(global_tmr_voter(2)(158));                                                             
 
                tmr_registers(0)(160)    <= not(global_tmr_voter(0)(159));                                                             
                tmr_registers(1)(160)    <= not(global_tmr_voter(1)(159));                                                             
                tmr_registers(2)(160)    <= not(global_tmr_voter(2)(159));                                                             
 
                tmr_registers(0)(161)    <= not(global_tmr_voter(0)(160));                                                             
                tmr_registers(1)(161)    <= not(global_tmr_voter(1)(160));                                                             
                tmr_registers(2)(161)    <= not(global_tmr_voter(2)(160));                                                             
 
                tmr_registers(0)(162)    <= not(global_tmr_voter(0)(161));                                                             
                tmr_registers(1)(162)    <= not(global_tmr_voter(1)(161));                                                             
                tmr_registers(2)(162)    <= not(global_tmr_voter(2)(161));                                                             
 
                tmr_registers(0)(163)    <= not(global_tmr_voter(0)(162));                                                             
                tmr_registers(1)(163)    <= not(global_tmr_voter(1)(162));                                                             
                tmr_registers(2)(163)    <= not(global_tmr_voter(2)(162));                                                             
 
                tmr_registers(0)(164)    <= not(global_tmr_voter(0)(163));                                                             
                tmr_registers(1)(164)    <= not(global_tmr_voter(1)(163));                                                             
                tmr_registers(2)(164)    <= not(global_tmr_voter(2)(163));                                                             
 
                tmr_registers(0)(165)    <= not(global_tmr_voter(0)(164));                                                             
                tmr_registers(1)(165)    <= not(global_tmr_voter(1)(164));                                                             
                tmr_registers(2)(165)    <= not(global_tmr_voter(2)(164));                                                             
 
                tmr_registers(0)(166)    <= not(global_tmr_voter(0)(165));                                                             
                tmr_registers(1)(166)    <= not(global_tmr_voter(1)(165));                                                             
                tmr_registers(2)(166)    <= not(global_tmr_voter(2)(165));                                                             
 
                tmr_registers(0)(167)    <= not(global_tmr_voter(0)(166));                                                             
                tmr_registers(1)(167)    <= not(global_tmr_voter(1)(166));                                                             
                tmr_registers(2)(167)    <= not(global_tmr_voter(2)(166));                                                             
 
                tmr_registers(0)(168)    <= not(global_tmr_voter(0)(167));                                                             
                tmr_registers(1)(168)    <= not(global_tmr_voter(1)(167));                                                             
                tmr_registers(2)(168)    <= not(global_tmr_voter(2)(167));                                                             
 
                tmr_registers(0)(169)    <= not(global_tmr_voter(0)(168));                                                             
                tmr_registers(1)(169)    <= not(global_tmr_voter(1)(168));                                                             
                tmr_registers(2)(169)    <= not(global_tmr_voter(2)(168));                                                             
 
                tmr_registers(0)(170)    <= not(global_tmr_voter(0)(169));                                                             
                tmr_registers(1)(170)    <= not(global_tmr_voter(1)(169));                                                             
                tmr_registers(2)(170)    <= not(global_tmr_voter(2)(169));                                                             
 
                tmr_registers(0)(171)    <= not(global_tmr_voter(0)(170));                                                             
                tmr_registers(1)(171)    <= not(global_tmr_voter(1)(170));                                                             
                tmr_registers(2)(171)    <= not(global_tmr_voter(2)(170));                                                             
 
                tmr_registers(0)(172)    <= not(global_tmr_voter(0)(171));                                                             
                tmr_registers(1)(172)    <= not(global_tmr_voter(1)(171));                                                             
                tmr_registers(2)(172)    <= not(global_tmr_voter(2)(171));                                                             
 
                tmr_registers(0)(173)    <= not(global_tmr_voter(0)(172));                                                             
                tmr_registers(1)(173)    <= not(global_tmr_voter(1)(172));                                                             
                tmr_registers(2)(173)    <= not(global_tmr_voter(2)(172));                                                             
 
                tmr_registers(0)(174)    <= not(global_tmr_voter(0)(173));                                                             
                tmr_registers(1)(174)    <= not(global_tmr_voter(1)(173));                                                             
                tmr_registers(2)(174)    <= not(global_tmr_voter(2)(173));                                                             
 
                tmr_registers(0)(175)    <= not(global_tmr_voter(0)(174));                                                             
                tmr_registers(1)(175)    <= not(global_tmr_voter(1)(174));                                                             
                tmr_registers(2)(175)    <= not(global_tmr_voter(2)(174));                                                             
 
                tmr_registers(0)(176)    <= not(global_tmr_voter(0)(175));                                                             
                tmr_registers(1)(176)    <= not(global_tmr_voter(1)(175));                                                             
                tmr_registers(2)(176)    <= not(global_tmr_voter(2)(175));                                                             
 
                tmr_registers(0)(177)    <= not(global_tmr_voter(0)(176));                                                             
                tmr_registers(1)(177)    <= not(global_tmr_voter(1)(176));                                                             
                tmr_registers(2)(177)    <= not(global_tmr_voter(2)(176));                                                             
 
                tmr_registers(0)(178)    <= not(global_tmr_voter(0)(177));                                                             
                tmr_registers(1)(178)    <= not(global_tmr_voter(1)(177));                                                             
                tmr_registers(2)(178)    <= not(global_tmr_voter(2)(177));                                                             
 
                tmr_registers(0)(179)    <= not(global_tmr_voter(0)(178));                                                             
                tmr_registers(1)(179)    <= not(global_tmr_voter(1)(178));                                                             
                tmr_registers(2)(179)    <= not(global_tmr_voter(2)(178));                                                             
 
                tmr_registers(0)(180)    <= not(global_tmr_voter(0)(179));                                                             
                tmr_registers(1)(180)    <= not(global_tmr_voter(1)(179));                                                             
                tmr_registers(2)(180)    <= not(global_tmr_voter(2)(179));                                                             
 
                tmr_registers(0)(181)    <= not(global_tmr_voter(0)(180));                                                             
                tmr_registers(1)(181)    <= not(global_tmr_voter(1)(180));                                                             
                tmr_registers(2)(181)    <= not(global_tmr_voter(2)(180));                                                             
 
                tmr_registers(0)(182)    <= not(global_tmr_voter(0)(181));                                                             
                tmr_registers(1)(182)    <= not(global_tmr_voter(1)(181));                                                             
                tmr_registers(2)(182)    <= not(global_tmr_voter(2)(181));                                                             
 
                tmr_registers(0)(183)    <= not(global_tmr_voter(0)(182));                                                             
                tmr_registers(1)(183)    <= not(global_tmr_voter(1)(182));                                                             
                tmr_registers(2)(183)    <= not(global_tmr_voter(2)(182));                                                             
 
                tmr_registers(0)(184)    <= not(global_tmr_voter(0)(183));                                                             
                tmr_registers(1)(184)    <= not(global_tmr_voter(1)(183));                                                             
                tmr_registers(2)(184)    <= not(global_tmr_voter(2)(183));                                                             
 
                tmr_registers(0)(185)    <= not(global_tmr_voter(0)(184));                                                             
                tmr_registers(1)(185)    <= not(global_tmr_voter(1)(184));                                                             
                tmr_registers(2)(185)    <= not(global_tmr_voter(2)(184));                                                             
 
                tmr_registers(0)(186)    <= not(global_tmr_voter(0)(185));                                                             
                tmr_registers(1)(186)    <= not(global_tmr_voter(1)(185));                                                             
                tmr_registers(2)(186)    <= not(global_tmr_voter(2)(185));                                                             
 
                tmr_registers(0)(187)    <= not(global_tmr_voter(0)(186));                                                             
                tmr_registers(1)(187)    <= not(global_tmr_voter(1)(186));                                                             
                tmr_registers(2)(187)    <= not(global_tmr_voter(2)(186));                                                             
 
                tmr_registers(0)(188)    <= not(global_tmr_voter(0)(187));                                                             
                tmr_registers(1)(188)    <= not(global_tmr_voter(1)(187));                                                             
                tmr_registers(2)(188)    <= not(global_tmr_voter(2)(187));                                                             
 
                tmr_registers(0)(189)    <= not(global_tmr_voter(0)(188));                                                             
                tmr_registers(1)(189)    <= not(global_tmr_voter(1)(188));                                                             
                tmr_registers(2)(189)    <= not(global_tmr_voter(2)(188));                                                             
 
                tmr_registers(0)(190)    <= not(global_tmr_voter(0)(189));                                                             
                tmr_registers(1)(190)    <= not(global_tmr_voter(1)(189));                                                             
                tmr_registers(2)(190)    <= not(global_tmr_voter(2)(189));                                                             
 
                tmr_registers(0)(191)    <= not(global_tmr_voter(0)(190));                                                             
                tmr_registers(1)(191)    <= not(global_tmr_voter(1)(190));                                                             
                tmr_registers(2)(191)    <= not(global_tmr_voter(2)(190));                                                             
 
                tmr_registers(0)(192)    <= not(global_tmr_voter(0)(191));                                                             
                tmr_registers(1)(192)    <= not(global_tmr_voter(1)(191));                                                             
                tmr_registers(2)(192)    <= not(global_tmr_voter(2)(191));                                                             
 
                tmr_registers(0)(193)    <= not(global_tmr_voter(0)(192));                                                             
                tmr_registers(1)(193)    <= not(global_tmr_voter(1)(192));                                                             
                tmr_registers(2)(193)    <= not(global_tmr_voter(2)(192));                                                             
 
                tmr_registers(0)(194)    <= not(global_tmr_voter(0)(193));                                                             
                tmr_registers(1)(194)    <= not(global_tmr_voter(1)(193));                                                             
                tmr_registers(2)(194)    <= not(global_tmr_voter(2)(193));                                                             
 
                tmr_registers(0)(195)    <= not(global_tmr_voter(0)(194));                                                             
                tmr_registers(1)(195)    <= not(global_tmr_voter(1)(194));                                                             
                tmr_registers(2)(195)    <= not(global_tmr_voter(2)(194));                                                             
 
                tmr_registers(0)(196)    <= not(global_tmr_voter(0)(195));                                                             
                tmr_registers(1)(196)    <= not(global_tmr_voter(1)(195));                                                             
                tmr_registers(2)(196)    <= not(global_tmr_voter(2)(195));                                                             
 
                tmr_registers(0)(197)    <= not(global_tmr_voter(0)(196));                                                             
                tmr_registers(1)(197)    <= not(global_tmr_voter(1)(196));                                                             
                tmr_registers(2)(197)    <= not(global_tmr_voter(2)(196));                                                             
 
                tmr_registers(0)(198)    <= not(global_tmr_voter(0)(197));                                                             
                tmr_registers(1)(198)    <= not(global_tmr_voter(1)(197));                                                             
                tmr_registers(2)(198)    <= not(global_tmr_voter(2)(197));                                                             
 
                tmr_registers(0)(199)    <= not(global_tmr_voter(0)(198));                                                             
                tmr_registers(1)(199)    <= not(global_tmr_voter(1)(198));                                                             
                tmr_registers(2)(199)    <= not(global_tmr_voter(2)(198));                                                             
 
                tmr_registers(0)(200)    <= not(global_tmr_voter(0)(199));                                                             
                tmr_registers(1)(200)    <= not(global_tmr_voter(1)(199));                                                             
                tmr_registers(2)(200)    <= not(global_tmr_voter(2)(199));                                                             
 
                tmr_registers(0)(201)    <= not(global_tmr_voter(0)(200));                                                             
                tmr_registers(1)(201)    <= not(global_tmr_voter(1)(200));                                                             
                tmr_registers(2)(201)    <= not(global_tmr_voter(2)(200));                                                             
 
                tmr_registers(0)(202)    <= not(global_tmr_voter(0)(201));                                                             
                tmr_registers(1)(202)    <= not(global_tmr_voter(1)(201));                                                             
                tmr_registers(2)(202)    <= not(global_tmr_voter(2)(201));                                                             
 
                tmr_registers(0)(203)    <= not(global_tmr_voter(0)(202));                                                             
                tmr_registers(1)(203)    <= not(global_tmr_voter(1)(202));                                                             
                tmr_registers(2)(203)    <= not(global_tmr_voter(2)(202));                                                             
 
                tmr_registers(0)(204)    <= not(global_tmr_voter(0)(203));                                                             
                tmr_registers(1)(204)    <= not(global_tmr_voter(1)(203));                                                             
                tmr_registers(2)(204)    <= not(global_tmr_voter(2)(203));                                                             
 
                tmr_registers(0)(205)    <= not(global_tmr_voter(0)(204));                                                             
                tmr_registers(1)(205)    <= not(global_tmr_voter(1)(204));                                                             
                tmr_registers(2)(205)    <= not(global_tmr_voter(2)(204));                                                             
 
                tmr_registers(0)(206)    <= not(global_tmr_voter(0)(205));                                                             
                tmr_registers(1)(206)    <= not(global_tmr_voter(1)(205));                                                             
                tmr_registers(2)(206)    <= not(global_tmr_voter(2)(205));                                                             
 
                tmr_registers(0)(207)    <= not(global_tmr_voter(0)(206));                                                             
                tmr_registers(1)(207)    <= not(global_tmr_voter(1)(206));                                                             
                tmr_registers(2)(207)    <= not(global_tmr_voter(2)(206));                                                             
 
                tmr_registers(0)(208)    <= not(global_tmr_voter(0)(207));                                                             
                tmr_registers(1)(208)    <= not(global_tmr_voter(1)(207));                                                             
                tmr_registers(2)(208)    <= not(global_tmr_voter(2)(207));                                                             
 
                tmr_registers(0)(209)    <= not(global_tmr_voter(0)(208));                                                             
                tmr_registers(1)(209)    <= not(global_tmr_voter(1)(208));                                                             
                tmr_registers(2)(209)    <= not(global_tmr_voter(2)(208));                                                             
 
                tmr_registers(0)(210)    <= not(global_tmr_voter(0)(209));                                                             
                tmr_registers(1)(210)    <= not(global_tmr_voter(1)(209));                                                             
                tmr_registers(2)(210)    <= not(global_tmr_voter(2)(209));                                                             
 
                tmr_registers(0)(211)    <= not(global_tmr_voter(0)(210));                                                             
                tmr_registers(1)(211)    <= not(global_tmr_voter(1)(210));                                                             
                tmr_registers(2)(211)    <= not(global_tmr_voter(2)(210));                                                             
 
                tmr_registers(0)(212)    <= not(global_tmr_voter(0)(211));                                                             
                tmr_registers(1)(212)    <= not(global_tmr_voter(1)(211));                                                             
                tmr_registers(2)(212)    <= not(global_tmr_voter(2)(211));                                                             
 
                tmr_registers(0)(213)    <= not(global_tmr_voter(0)(212));                                                             
                tmr_registers(1)(213)    <= not(global_tmr_voter(1)(212));                                                             
                tmr_registers(2)(213)    <= not(global_tmr_voter(2)(212));                                                             
 
                tmr_registers(0)(214)    <= not(global_tmr_voter(0)(213));                                                             
                tmr_registers(1)(214)    <= not(global_tmr_voter(1)(213));                                                             
                tmr_registers(2)(214)    <= not(global_tmr_voter(2)(213));                                                             
 
                tmr_registers(0)(215)    <= not(global_tmr_voter(0)(214));                                                             
                tmr_registers(1)(215)    <= not(global_tmr_voter(1)(214));                                                             
                tmr_registers(2)(215)    <= not(global_tmr_voter(2)(214));                                                             
 
                tmr_registers(0)(216)    <= not(global_tmr_voter(0)(215));                                                             
                tmr_registers(1)(216)    <= not(global_tmr_voter(1)(215));                                                             
                tmr_registers(2)(216)    <= not(global_tmr_voter(2)(215));                                                             
 
                tmr_registers(0)(217)    <= not(global_tmr_voter(0)(216));                                                             
                tmr_registers(1)(217)    <= not(global_tmr_voter(1)(216));                                                             
                tmr_registers(2)(217)    <= not(global_tmr_voter(2)(216));                                                             
 
                tmr_registers(0)(218)    <= not(global_tmr_voter(0)(217));                                                             
                tmr_registers(1)(218)    <= not(global_tmr_voter(1)(217));                                                             
                tmr_registers(2)(218)    <= not(global_tmr_voter(2)(217));                                                             
 
                tmr_registers(0)(219)    <= not(global_tmr_voter(0)(218));                                                             
                tmr_registers(1)(219)    <= not(global_tmr_voter(1)(218));                                                             
                tmr_registers(2)(219)    <= not(global_tmr_voter(2)(218));                                                             
 
                tmr_registers(0)(220)    <= not(global_tmr_voter(0)(219));                                                             
                tmr_registers(1)(220)    <= not(global_tmr_voter(1)(219));                                                             
                tmr_registers(2)(220)    <= not(global_tmr_voter(2)(219));                                                             
 
                tmr_registers(0)(221)    <= not(global_tmr_voter(0)(220));                                                             
                tmr_registers(1)(221)    <= not(global_tmr_voter(1)(220));                                                             
                tmr_registers(2)(221)    <= not(global_tmr_voter(2)(220));                                                             
 
                tmr_registers(0)(222)    <= not(global_tmr_voter(0)(221));                                                             
                tmr_registers(1)(222)    <= not(global_tmr_voter(1)(221));                                                             
                tmr_registers(2)(222)    <= not(global_tmr_voter(2)(221));                                                             
 
                tmr_registers(0)(223)    <= not(global_tmr_voter(0)(222));                                                             
                tmr_registers(1)(223)    <= not(global_tmr_voter(1)(222));                                                             
                tmr_registers(2)(223)    <= not(global_tmr_voter(2)(222));                                                             
 
                tmr_registers(0)(224)    <= not(global_tmr_voter(0)(223));                                                             
                tmr_registers(1)(224)    <= not(global_tmr_voter(1)(223));                                                             
                tmr_registers(2)(224)    <= not(global_tmr_voter(2)(223));                                                             
 
                tmr_registers(0)(225)    <= not(global_tmr_voter(0)(224));                                                             
                tmr_registers(1)(225)    <= not(global_tmr_voter(1)(224));                                                             
                tmr_registers(2)(225)    <= not(global_tmr_voter(2)(224));                                                             
 
                tmr_registers(0)(226)    <= not(global_tmr_voter(0)(225));                                                             
                tmr_registers(1)(226)    <= not(global_tmr_voter(1)(225));                                                             
                tmr_registers(2)(226)    <= not(global_tmr_voter(2)(225));                                                             
 
                tmr_registers(0)(227)    <= not(global_tmr_voter(0)(226));                                                             
                tmr_registers(1)(227)    <= not(global_tmr_voter(1)(226));                                                             
                tmr_registers(2)(227)    <= not(global_tmr_voter(2)(226));                                                             
 
                tmr_registers(0)(228)    <= not(global_tmr_voter(0)(227));                                                             
                tmr_registers(1)(228)    <= not(global_tmr_voter(1)(227));                                                             
                tmr_registers(2)(228)    <= not(global_tmr_voter(2)(227));                                                             
 
                tmr_registers(0)(229)    <= not(global_tmr_voter(0)(228));                                                             
                tmr_registers(1)(229)    <= not(global_tmr_voter(1)(228));                                                             
                tmr_registers(2)(229)    <= not(global_tmr_voter(2)(228));                                                             
 
                tmr_registers(0)(230)    <= not(global_tmr_voter(0)(229));                                                             
                tmr_registers(1)(230)    <= not(global_tmr_voter(1)(229));                                                             
                tmr_registers(2)(230)    <= not(global_tmr_voter(2)(229));                                                             
 
                tmr_registers(0)(231)    <= not(global_tmr_voter(0)(230));                                                             
                tmr_registers(1)(231)    <= not(global_tmr_voter(1)(230));                                                             
                tmr_registers(2)(231)    <= not(global_tmr_voter(2)(230));                                                             
 
                tmr_registers(0)(232)    <= not(global_tmr_voter(0)(231));                                                             
                tmr_registers(1)(232)    <= not(global_tmr_voter(1)(231));                                                             
                tmr_registers(2)(232)    <= not(global_tmr_voter(2)(231));                                                             
 
                tmr_registers(0)(233)    <= not(global_tmr_voter(0)(232));                                                             
                tmr_registers(1)(233)    <= not(global_tmr_voter(1)(232));                                                             
                tmr_registers(2)(233)    <= not(global_tmr_voter(2)(232));                                                             
 
                tmr_registers(0)(234)    <= not(global_tmr_voter(0)(233));                                                             
                tmr_registers(1)(234)    <= not(global_tmr_voter(1)(233));                                                             
                tmr_registers(2)(234)    <= not(global_tmr_voter(2)(233));                                                             
 
                tmr_registers(0)(235)    <= not(global_tmr_voter(0)(234));                                                             
                tmr_registers(1)(235)    <= not(global_tmr_voter(1)(234));                                                             
                tmr_registers(2)(235)    <= not(global_tmr_voter(2)(234));                                                             
 
                tmr_registers(0)(236)    <= not(global_tmr_voter(0)(235));                                                             
                tmr_registers(1)(236)    <= not(global_tmr_voter(1)(235));                                                             
                tmr_registers(2)(236)    <= not(global_tmr_voter(2)(235));                                                             
 
                tmr_registers(0)(237)    <= not(global_tmr_voter(0)(236));                                                             
                tmr_registers(1)(237)    <= not(global_tmr_voter(1)(236));                                                             
                tmr_registers(2)(237)    <= not(global_tmr_voter(2)(236));                                                             
 
                tmr_registers(0)(238)    <= not(global_tmr_voter(0)(237));                                                             
                tmr_registers(1)(238)    <= not(global_tmr_voter(1)(237));                                                             
                tmr_registers(2)(238)    <= not(global_tmr_voter(2)(237));                                                             
 
                tmr_registers(0)(239)    <= not(global_tmr_voter(0)(238));                                                             
                tmr_registers(1)(239)    <= not(global_tmr_voter(1)(238));                                                             
                tmr_registers(2)(239)    <= not(global_tmr_voter(2)(238));                                                             
 
                tmr_registers(0)(240)    <= not(global_tmr_voter(0)(239));                                                             
                tmr_registers(1)(240)    <= not(global_tmr_voter(1)(239));                                                             
                tmr_registers(2)(240)    <= not(global_tmr_voter(2)(239));                                                             
 
                tmr_registers(0)(241)    <= not(global_tmr_voter(0)(240));                                                             
                tmr_registers(1)(241)    <= not(global_tmr_voter(1)(240));                                                             
                tmr_registers(2)(241)    <= not(global_tmr_voter(2)(240));                                                             
 
                tmr_registers(0)(242)    <= not(global_tmr_voter(0)(241));                                                             
                tmr_registers(1)(242)    <= not(global_tmr_voter(1)(241));                                                             
                tmr_registers(2)(242)    <= not(global_tmr_voter(2)(241));                                                             
 
                tmr_registers(0)(243)    <= not(global_tmr_voter(0)(242));                                                             
                tmr_registers(1)(243)    <= not(global_tmr_voter(1)(242));                                                             
                tmr_registers(2)(243)    <= not(global_tmr_voter(2)(242));                                                             
 
                tmr_registers(0)(244)    <= not(global_tmr_voter(0)(243));                                                             
                tmr_registers(1)(244)    <= not(global_tmr_voter(1)(243));                                                             
                tmr_registers(2)(244)    <= not(global_tmr_voter(2)(243));                                                             
 
                tmr_registers(0)(245)    <= not(global_tmr_voter(0)(244));                                                             
                tmr_registers(1)(245)    <= not(global_tmr_voter(1)(244));                                                             
                tmr_registers(2)(245)    <= not(global_tmr_voter(2)(244));                                                             
 
                tmr_registers(0)(246)    <= not(global_tmr_voter(0)(245));                                                             
                tmr_registers(1)(246)    <= not(global_tmr_voter(1)(245));                                                             
                tmr_registers(2)(246)    <= not(global_tmr_voter(2)(245));                                                             
 
                tmr_registers(0)(247)    <= not(global_tmr_voter(0)(246));                                                             
                tmr_registers(1)(247)    <= not(global_tmr_voter(1)(246));                                                             
                tmr_registers(2)(247)    <= not(global_tmr_voter(2)(246));                                                             
 
                tmr_registers(0)(248)    <= not(global_tmr_voter(0)(247));                                                             
                tmr_registers(1)(248)    <= not(global_tmr_voter(1)(247));                                                             
                tmr_registers(2)(248)    <= not(global_tmr_voter(2)(247));                                                             
 
                tmr_registers(0)(249)    <= not(global_tmr_voter(0)(248));                                                             
                tmr_registers(1)(249)    <= not(global_tmr_voter(1)(248));                                                             
                tmr_registers(2)(249)    <= not(global_tmr_voter(2)(248));                                                             
 
                tmr_registers(0)(250)    <= not(global_tmr_voter(0)(249));                                                             
                tmr_registers(1)(250)    <= not(global_tmr_voter(1)(249));                                                             
                tmr_registers(2)(250)    <= not(global_tmr_voter(2)(249));                                                             
 
                tmr_registers(0)(251)    <= not(global_tmr_voter(0)(250));                                                             
                tmr_registers(1)(251)    <= not(global_tmr_voter(1)(250));                                                             
                tmr_registers(2)(251)    <= not(global_tmr_voter(2)(250));                                                             
 
                tmr_registers(0)(252)    <= not(global_tmr_voter(0)(251));                                                             
                tmr_registers(1)(252)    <= not(global_tmr_voter(1)(251));                                                             
                tmr_registers(2)(252)    <= not(global_tmr_voter(2)(251));                                                             
 
                tmr_registers(0)(253)    <= not(global_tmr_voter(0)(252));                                                             
                tmr_registers(1)(253)    <= not(global_tmr_voter(1)(252));                                                             
                tmr_registers(2)(253)    <= not(global_tmr_voter(2)(252));                                                             
 
                tmr_registers(0)(254)    <= not(global_tmr_voter(0)(253));                                                             
                tmr_registers(1)(254)    <= not(global_tmr_voter(1)(253));                                                             
                tmr_registers(2)(254)    <= not(global_tmr_voter(2)(253));                                                             
 
                tmr_registers(0)(255)    <= not(global_tmr_voter(0)(254));                                                             
                tmr_registers(1)(255)    <= not(global_tmr_voter(1)(254));                                                             
                tmr_registers(2)(255)    <= not(global_tmr_voter(2)(254));                                                             
 
                tmr_registers(0)(256)    <= not(global_tmr_voter(0)(255));                                                             
                tmr_registers(1)(256)    <= not(global_tmr_voter(1)(255));                                                             
                tmr_registers(2)(256)    <= not(global_tmr_voter(2)(255));                                                             
 
                tmr_registers(0)(257)    <= not(global_tmr_voter(0)(256));                                                             
                tmr_registers(1)(257)    <= not(global_tmr_voter(1)(256));                                                             
                tmr_registers(2)(257)    <= not(global_tmr_voter(2)(256));                                                             
 
                tmr_registers(0)(258)    <= not(global_tmr_voter(0)(257));                                                             
                tmr_registers(1)(258)    <= not(global_tmr_voter(1)(257));                                                             
                tmr_registers(2)(258)    <= not(global_tmr_voter(2)(257));                                                             
 
                tmr_registers(0)(259)    <= not(global_tmr_voter(0)(258));                                                             
                tmr_registers(1)(259)    <= not(global_tmr_voter(1)(258));                                                             
                tmr_registers(2)(259)    <= not(global_tmr_voter(2)(258));                                                             
 
                tmr_registers(0)(260)    <= not(global_tmr_voter(0)(259));                                                             
                tmr_registers(1)(260)    <= not(global_tmr_voter(1)(259));                                                             
                tmr_registers(2)(260)    <= not(global_tmr_voter(2)(259));                                                             
 
                tmr_registers(0)(261)    <= not(global_tmr_voter(0)(260));                                                             
                tmr_registers(1)(261)    <= not(global_tmr_voter(1)(260));                                                             
                tmr_registers(2)(261)    <= not(global_tmr_voter(2)(260));                                                             
 
                tmr_registers(0)(262)    <= not(global_tmr_voter(0)(261));                                                             
                tmr_registers(1)(262)    <= not(global_tmr_voter(1)(261));                                                             
                tmr_registers(2)(262)    <= not(global_tmr_voter(2)(261));                                                             
 
                tmr_registers(0)(263)    <= not(global_tmr_voter(0)(262));                                                             
                tmr_registers(1)(263)    <= not(global_tmr_voter(1)(262));                                                             
                tmr_registers(2)(263)    <= not(global_tmr_voter(2)(262));                                                             
 
                tmr_registers(0)(264)    <= not(global_tmr_voter(0)(263));                                                             
                tmr_registers(1)(264)    <= not(global_tmr_voter(1)(263));                                                             
                tmr_registers(2)(264)    <= not(global_tmr_voter(2)(263));                                                             
 
                tmr_registers(0)(265)    <= not(global_tmr_voter(0)(264));                                                             
                tmr_registers(1)(265)    <= not(global_tmr_voter(1)(264));                                                             
                tmr_registers(2)(265)    <= not(global_tmr_voter(2)(264));                                                             
 
                tmr_registers(0)(266)    <= not(global_tmr_voter(0)(265));                                                             
                tmr_registers(1)(266)    <= not(global_tmr_voter(1)(265));                                                             
                tmr_registers(2)(266)    <= not(global_tmr_voter(2)(265));                                                             
 
                tmr_registers(0)(267)    <= not(global_tmr_voter(0)(266));                                                             
                tmr_registers(1)(267)    <= not(global_tmr_voter(1)(266));                                                             
                tmr_registers(2)(267)    <= not(global_tmr_voter(2)(266));                                                             
 
                tmr_registers(0)(268)    <= not(global_tmr_voter(0)(267));                                                             
                tmr_registers(1)(268)    <= not(global_tmr_voter(1)(267));                                                             
                tmr_registers(2)(268)    <= not(global_tmr_voter(2)(267));                                                             
 
                tmr_registers(0)(269)    <= not(global_tmr_voter(0)(268));                                                             
                tmr_registers(1)(269)    <= not(global_tmr_voter(1)(268));                                                             
                tmr_registers(2)(269)    <= not(global_tmr_voter(2)(268));                                                             
 
                tmr_registers(0)(270)    <= not(global_tmr_voter(0)(269));                                                             
                tmr_registers(1)(270)    <= not(global_tmr_voter(1)(269));                                                             
                tmr_registers(2)(270)    <= not(global_tmr_voter(2)(269));                                                             
 
                tmr_registers(0)(271)    <= not(global_tmr_voter(0)(270));                                                             
                tmr_registers(1)(271)    <= not(global_tmr_voter(1)(270));                                                             
                tmr_registers(2)(271)    <= not(global_tmr_voter(2)(270));                                                             
 
                tmr_registers(0)(272)    <= not(global_tmr_voter(0)(271));                                                             
                tmr_registers(1)(272)    <= not(global_tmr_voter(1)(271));                                                             
                tmr_registers(2)(272)    <= not(global_tmr_voter(2)(271));                                                             
 
                tmr_registers(0)(273)    <= not(global_tmr_voter(0)(272));                                                             
                tmr_registers(1)(273)    <= not(global_tmr_voter(1)(272));                                                             
                tmr_registers(2)(273)    <= not(global_tmr_voter(2)(272));                                                             
 
                tmr_registers(0)(274)    <= not(global_tmr_voter(0)(273));                                                             
                tmr_registers(1)(274)    <= not(global_tmr_voter(1)(273));                                                             
                tmr_registers(2)(274)    <= not(global_tmr_voter(2)(273));                                                             
 
                tmr_registers(0)(275)    <= not(global_tmr_voter(0)(274));                                                             
                tmr_registers(1)(275)    <= not(global_tmr_voter(1)(274));                                                             
                tmr_registers(2)(275)    <= not(global_tmr_voter(2)(274));                                                             
 
                tmr_registers(0)(276)    <= not(global_tmr_voter(0)(275));                                                             
                tmr_registers(1)(276)    <= not(global_tmr_voter(1)(275));                                                             
                tmr_registers(2)(276)    <= not(global_tmr_voter(2)(275));                                                             
 
                tmr_registers(0)(277)    <= not(global_tmr_voter(0)(276));                                                             
                tmr_registers(1)(277)    <= not(global_tmr_voter(1)(276));                                                             
                tmr_registers(2)(277)    <= not(global_tmr_voter(2)(276));                                                             
 
                tmr_registers(0)(278)    <= not(global_tmr_voter(0)(277));                                                             
                tmr_registers(1)(278)    <= not(global_tmr_voter(1)(277));                                                             
                tmr_registers(2)(278)    <= not(global_tmr_voter(2)(277));                                                             
 
                tmr_registers(0)(279)    <= not(global_tmr_voter(0)(278));                                                             
                tmr_registers(1)(279)    <= not(global_tmr_voter(1)(278));                                                             
                tmr_registers(2)(279)    <= not(global_tmr_voter(2)(278));                                                             
 
                tmr_registers(0)(280)    <= not(global_tmr_voter(0)(279));                                                             
                tmr_registers(1)(280)    <= not(global_tmr_voter(1)(279));                                                             
                tmr_registers(2)(280)    <= not(global_tmr_voter(2)(279));                                                             
 
                tmr_registers(0)(281)    <= not(global_tmr_voter(0)(280));                                                             
                tmr_registers(1)(281)    <= not(global_tmr_voter(1)(280));                                                             
                tmr_registers(2)(281)    <= not(global_tmr_voter(2)(280));                                                             
 
                tmr_registers(0)(282)    <= not(global_tmr_voter(0)(281));                                                             
                tmr_registers(1)(282)    <= not(global_tmr_voter(1)(281));                                                             
                tmr_registers(2)(282)    <= not(global_tmr_voter(2)(281));                                                             
 
                tmr_registers(0)(283)    <= not(global_tmr_voter(0)(282));                                                             
                tmr_registers(1)(283)    <= not(global_tmr_voter(1)(282));                                                             
                tmr_registers(2)(283)    <= not(global_tmr_voter(2)(282));                                                             
 
                tmr_registers(0)(284)    <= not(global_tmr_voter(0)(283));                                                             
                tmr_registers(1)(284)    <= not(global_tmr_voter(1)(283));                                                             
                tmr_registers(2)(284)    <= not(global_tmr_voter(2)(283));                                                             
 
                tmr_registers(0)(285)    <= not(global_tmr_voter(0)(284));                                                             
                tmr_registers(1)(285)    <= not(global_tmr_voter(1)(284));                                                             
                tmr_registers(2)(285)    <= not(global_tmr_voter(2)(284));                                                             
 
                tmr_registers(0)(286)    <= not(global_tmr_voter(0)(285));                                                             
                tmr_registers(1)(286)    <= not(global_tmr_voter(1)(285));                                                             
                tmr_registers(2)(286)    <= not(global_tmr_voter(2)(285));                                                             
 
                tmr_registers(0)(287)    <= not(global_tmr_voter(0)(286));                                                             
                tmr_registers(1)(287)    <= not(global_tmr_voter(1)(286));                                                             
                tmr_registers(2)(287)    <= not(global_tmr_voter(2)(286));                                                             
 
                tmr_registers(0)(288)    <= not(global_tmr_voter(0)(287));                                                             
                tmr_registers(1)(288)    <= not(global_tmr_voter(1)(287));                                                             
                tmr_registers(2)(288)    <= not(global_tmr_voter(2)(287));                                                             
 
                tmr_registers(0)(289)    <= not(global_tmr_voter(0)(288));                                                             
                tmr_registers(1)(289)    <= not(global_tmr_voter(1)(288));                                                             
                tmr_registers(2)(289)    <= not(global_tmr_voter(2)(288));                                                             
 
                tmr_registers(0)(290)    <= not(global_tmr_voter(0)(289));                                                             
                tmr_registers(1)(290)    <= not(global_tmr_voter(1)(289));                                                             
                tmr_registers(2)(290)    <= not(global_tmr_voter(2)(289));                                                             
 
                tmr_registers(0)(291)    <= not(global_tmr_voter(0)(290));                                                             
                tmr_registers(1)(291)    <= not(global_tmr_voter(1)(290));                                                             
                tmr_registers(2)(291)    <= not(global_tmr_voter(2)(290));                                                             
 
                tmr_registers(0)(292)    <= not(global_tmr_voter(0)(291));                                                             
                tmr_registers(1)(292)    <= not(global_tmr_voter(1)(291));                                                             
                tmr_registers(2)(292)    <= not(global_tmr_voter(2)(291));                                                             
 
                tmr_registers(0)(293)    <= not(global_tmr_voter(0)(292));                                                             
                tmr_registers(1)(293)    <= not(global_tmr_voter(1)(292));                                                             
                tmr_registers(2)(293)    <= not(global_tmr_voter(2)(292));                                                             
 
                tmr_registers(0)(294)    <= not(global_tmr_voter(0)(293));                                                             
                tmr_registers(1)(294)    <= not(global_tmr_voter(1)(293));                                                             
                tmr_registers(2)(294)    <= not(global_tmr_voter(2)(293));                                                             
 
                tmr_registers(0)(295)    <= not(global_tmr_voter(0)(294));                                                             
                tmr_registers(1)(295)    <= not(global_tmr_voter(1)(294));                                                             
                tmr_registers(2)(295)    <= not(global_tmr_voter(2)(294));                                                             
 
                tmr_registers(0)(296)    <= not(global_tmr_voter(0)(295));                                                             
                tmr_registers(1)(296)    <= not(global_tmr_voter(1)(295));                                                             
                tmr_registers(2)(296)    <= not(global_tmr_voter(2)(295));                                                             
 
                tmr_registers(0)(297)    <= not(global_tmr_voter(0)(296));                                                             
                tmr_registers(1)(297)    <= not(global_tmr_voter(1)(296));                                                             
                tmr_registers(2)(297)    <= not(global_tmr_voter(2)(296));                                                             
 
                tmr_registers(0)(298)    <= not(global_tmr_voter(0)(297));                                                             
                tmr_registers(1)(298)    <= not(global_tmr_voter(1)(297));                                                             
                tmr_registers(2)(298)    <= not(global_tmr_voter(2)(297));                                                             
 
                tmr_registers(0)(299)    <= not(global_tmr_voter(0)(298));                                                             
                tmr_registers(1)(299)    <= not(global_tmr_voter(1)(298));                                                             
                tmr_registers(2)(299)    <= not(global_tmr_voter(2)(298));                                                             
 
                tmr_registers(0)(300)    <= not(global_tmr_voter(0)(299));                                                             
                tmr_registers(1)(300)    <= not(global_tmr_voter(1)(299));                                                             
                tmr_registers(2)(300)    <= not(global_tmr_voter(2)(299));                                                             
 
                tmr_registers(0)(301)    <= not(global_tmr_voter(0)(300));                                                             
                tmr_registers(1)(301)    <= not(global_tmr_voter(1)(300));                                                             
                tmr_registers(2)(301)    <= not(global_tmr_voter(2)(300));                                                             
 
                tmr_registers(0)(302)    <= not(global_tmr_voter(0)(301));                                                             
                tmr_registers(1)(302)    <= not(global_tmr_voter(1)(301));                                                             
                tmr_registers(2)(302)    <= not(global_tmr_voter(2)(301));                                                             
 
                tmr_registers(0)(303)    <= not(global_tmr_voter(0)(302));                                                             
                tmr_registers(1)(303)    <= not(global_tmr_voter(1)(302));                                                             
                tmr_registers(2)(303)    <= not(global_tmr_voter(2)(302));                                                             
 
                tmr_registers(0)(304)    <= not(global_tmr_voter(0)(303));                                                             
                tmr_registers(1)(304)    <= not(global_tmr_voter(1)(303));                                                             
                tmr_registers(2)(304)    <= not(global_tmr_voter(2)(303));                                                             
 
                tmr_registers(0)(305)    <= not(global_tmr_voter(0)(304));                                                             
                tmr_registers(1)(305)    <= not(global_tmr_voter(1)(304));                                                             
                tmr_registers(2)(305)    <= not(global_tmr_voter(2)(304));                                                             
 
                tmr_registers(0)(306)    <= not(global_tmr_voter(0)(305));                                                             
                tmr_registers(1)(306)    <= not(global_tmr_voter(1)(305));                                                             
                tmr_registers(2)(306)    <= not(global_tmr_voter(2)(305));                                                             
 
                tmr_registers(0)(307)    <= not(global_tmr_voter(0)(306));                                                             
                tmr_registers(1)(307)    <= not(global_tmr_voter(1)(306));                                                             
                tmr_registers(2)(307)    <= not(global_tmr_voter(2)(306));                                                             
 
                tmr_registers(0)(308)    <= not(global_tmr_voter(0)(307));                                                             
                tmr_registers(1)(308)    <= not(global_tmr_voter(1)(307));                                                             
                tmr_registers(2)(308)    <= not(global_tmr_voter(2)(307));                                                             
 
                tmr_registers(0)(309)    <= not(global_tmr_voter(0)(308));                                                             
                tmr_registers(1)(309)    <= not(global_tmr_voter(1)(308));                                                             
                tmr_registers(2)(309)    <= not(global_tmr_voter(2)(308));                                                             
 
                tmr_registers(0)(310)    <= not(global_tmr_voter(0)(309));                                                             
                tmr_registers(1)(310)    <= not(global_tmr_voter(1)(309));                                                             
                tmr_registers(2)(310)    <= not(global_tmr_voter(2)(309));                                                             
 
                tmr_registers(0)(311)    <= not(global_tmr_voter(0)(310));                                                             
                tmr_registers(1)(311)    <= not(global_tmr_voter(1)(310));                                                             
                tmr_registers(2)(311)    <= not(global_tmr_voter(2)(310));                                                             
 
                tmr_registers(0)(312)    <= not(global_tmr_voter(0)(311));                                                             
                tmr_registers(1)(312)    <= not(global_tmr_voter(1)(311));                                                             
                tmr_registers(2)(312)    <= not(global_tmr_voter(2)(311));                                                             
 
                tmr_registers(0)(313)    <= not(global_tmr_voter(0)(312));                                                             
                tmr_registers(1)(313)    <= not(global_tmr_voter(1)(312));                                                             
                tmr_registers(2)(313)    <= not(global_tmr_voter(2)(312));                                                             
 
                tmr_registers(0)(314)    <= not(global_tmr_voter(0)(313));                                                             
                tmr_registers(1)(314)    <= not(global_tmr_voter(1)(313));                                                             
                tmr_registers(2)(314)    <= not(global_tmr_voter(2)(313));                                                             
 
                tmr_registers(0)(315)    <= not(global_tmr_voter(0)(314));                                                             
                tmr_registers(1)(315)    <= not(global_tmr_voter(1)(314));                                                             
                tmr_registers(2)(315)    <= not(global_tmr_voter(2)(314));                                                             
 
                tmr_registers(0)(316)    <= not(global_tmr_voter(0)(315));                                                             
                tmr_registers(1)(316)    <= not(global_tmr_voter(1)(315));                                                             
                tmr_registers(2)(316)    <= not(global_tmr_voter(2)(315));                                                             
 
                tmr_registers(0)(317)    <= not(global_tmr_voter(0)(316));                                                             
                tmr_registers(1)(317)    <= not(global_tmr_voter(1)(316));                                                             
                tmr_registers(2)(317)    <= not(global_tmr_voter(2)(316));                                                             
 
                tmr_registers(0)(318)    <= not(global_tmr_voter(0)(317));                                                             
                tmr_registers(1)(318)    <= not(global_tmr_voter(1)(317));                                                             
                tmr_registers(2)(318)    <= not(global_tmr_voter(2)(317));                                                             
 
                tmr_registers(0)(319)    <= not(global_tmr_voter(0)(318));                                                             
                tmr_registers(1)(319)    <= not(global_tmr_voter(1)(318));                                                             
                tmr_registers(2)(319)    <= not(global_tmr_voter(2)(318));                                                             
 
                tmr_registers(0)(320)    <= not(global_tmr_voter(0)(319));                                                             
                tmr_registers(1)(320)    <= not(global_tmr_voter(1)(319));                                                             
                tmr_registers(2)(320)    <= not(global_tmr_voter(2)(319));                                                             
 
                tmr_registers(0)(321)    <= not(global_tmr_voter(0)(320));                                                             
                tmr_registers(1)(321)    <= not(global_tmr_voter(1)(320));                                                             
                tmr_registers(2)(321)    <= not(global_tmr_voter(2)(320));                                                             
 
                tmr_registers(0)(322)    <= not(global_tmr_voter(0)(321));                                                             
                tmr_registers(1)(322)    <= not(global_tmr_voter(1)(321));                                                             
                tmr_registers(2)(322)    <= not(global_tmr_voter(2)(321));                                                             
 
                tmr_registers(0)(323)    <= not(global_tmr_voter(0)(322));                                                             
                tmr_registers(1)(323)    <= not(global_tmr_voter(1)(322));                                                             
                tmr_registers(2)(323)    <= not(global_tmr_voter(2)(322));                                                             
 
                tmr_registers(0)(324)    <= not(global_tmr_voter(0)(323));                                                             
                tmr_registers(1)(324)    <= not(global_tmr_voter(1)(323));                                                             
                tmr_registers(2)(324)    <= not(global_tmr_voter(2)(323));                                                             
 
                tmr_registers(0)(325)    <= not(global_tmr_voter(0)(324));                                                             
                tmr_registers(1)(325)    <= not(global_tmr_voter(1)(324));                                                             
                tmr_registers(2)(325)    <= not(global_tmr_voter(2)(324));                                                             
 
                tmr_registers(0)(326)    <= not(global_tmr_voter(0)(325));                                                             
                tmr_registers(1)(326)    <= not(global_tmr_voter(1)(325));                                                             
                tmr_registers(2)(326)    <= not(global_tmr_voter(2)(325));                                                             
 
                tmr_registers(0)(327)    <= not(global_tmr_voter(0)(326));                                                             
                tmr_registers(1)(327)    <= not(global_tmr_voter(1)(326));                                                             
                tmr_registers(2)(327)    <= not(global_tmr_voter(2)(326));                                                             
 
                tmr_registers(0)(328)    <= not(global_tmr_voter(0)(327));                                                             
                tmr_registers(1)(328)    <= not(global_tmr_voter(1)(327));                                                             
                tmr_registers(2)(328)    <= not(global_tmr_voter(2)(327));                                                             
 
                tmr_registers(0)(329)    <= not(global_tmr_voter(0)(328));                                                             
                tmr_registers(1)(329)    <= not(global_tmr_voter(1)(328));                                                             
                tmr_registers(2)(329)    <= not(global_tmr_voter(2)(328));                                                             
 
                tmr_registers(0)(330)    <= not(global_tmr_voter(0)(329));                                                             
                tmr_registers(1)(330)    <= not(global_tmr_voter(1)(329));                                                             
                tmr_registers(2)(330)    <= not(global_tmr_voter(2)(329));                                                             
 
                tmr_registers(0)(331)    <= not(global_tmr_voter(0)(330));                                                             
                tmr_registers(1)(331)    <= not(global_tmr_voter(1)(330));                                                             
                tmr_registers(2)(331)    <= not(global_tmr_voter(2)(330));                                                             
 
                tmr_registers(0)(332)    <= not(global_tmr_voter(0)(331));                                                             
                tmr_registers(1)(332)    <= not(global_tmr_voter(1)(331));                                                             
                tmr_registers(2)(332)    <= not(global_tmr_voter(2)(331));                                                             
 
                tmr_registers(0)(333)    <= not(global_tmr_voter(0)(332));                                                             
                tmr_registers(1)(333)    <= not(global_tmr_voter(1)(332));                                                             
                tmr_registers(2)(333)    <= not(global_tmr_voter(2)(332));                                                             
 
                tmr_registers(0)(334)    <= not(global_tmr_voter(0)(333));                                                             
                tmr_registers(1)(334)    <= not(global_tmr_voter(1)(333));                                                             
                tmr_registers(2)(334)    <= not(global_tmr_voter(2)(333));                                                             
 
                tmr_registers(0)(335)    <= not(global_tmr_voter(0)(334));                                                             
                tmr_registers(1)(335)    <= not(global_tmr_voter(1)(334));                                                             
                tmr_registers(2)(335)    <= not(global_tmr_voter(2)(334));                                                             
 
                tmr_registers(0)(336)    <= not(global_tmr_voter(0)(335));                                                             
                tmr_registers(1)(336)    <= not(global_tmr_voter(1)(335));                                                             
                tmr_registers(2)(336)    <= not(global_tmr_voter(2)(335));                                                             
 
                tmr_registers(0)(337)    <= not(global_tmr_voter(0)(336));                                                             
                tmr_registers(1)(337)    <= not(global_tmr_voter(1)(336));                                                             
                tmr_registers(2)(337)    <= not(global_tmr_voter(2)(336));                                                             
 
                tmr_registers(0)(338)    <= not(global_tmr_voter(0)(337));                                                             
                tmr_registers(1)(338)    <= not(global_tmr_voter(1)(337));                                                             
                tmr_registers(2)(338)    <= not(global_tmr_voter(2)(337));                                                             
 
                tmr_registers(0)(339)    <= not(global_tmr_voter(0)(338));                                                             
                tmr_registers(1)(339)    <= not(global_tmr_voter(1)(338));                                                             
                tmr_registers(2)(339)    <= not(global_tmr_voter(2)(338));                                                             
 
                tmr_registers(0)(340)    <= not(global_tmr_voter(0)(339));                                                             
                tmr_registers(1)(340)    <= not(global_tmr_voter(1)(339));                                                             
                tmr_registers(2)(340)    <= not(global_tmr_voter(2)(339));                                                             
 
                tmr_registers(0)(341)    <= not(global_tmr_voter(0)(340));                                                             
                tmr_registers(1)(341)    <= not(global_tmr_voter(1)(340));                                                             
                tmr_registers(2)(341)    <= not(global_tmr_voter(2)(340));                                                             
 
                tmr_registers(0)(342)    <= not(global_tmr_voter(0)(341));                                                             
                tmr_registers(1)(342)    <= not(global_tmr_voter(1)(341));                                                             
                tmr_registers(2)(342)    <= not(global_tmr_voter(2)(341));                                                             
 
                tmr_registers(0)(343)    <= not(global_tmr_voter(0)(342));                                                             
                tmr_registers(1)(343)    <= not(global_tmr_voter(1)(342));                                                             
                tmr_registers(2)(343)    <= not(global_tmr_voter(2)(342));                                                             
 
                tmr_registers(0)(344)    <= not(global_tmr_voter(0)(343));                                                             
                tmr_registers(1)(344)    <= not(global_tmr_voter(1)(343));                                                             
                tmr_registers(2)(344)    <= not(global_tmr_voter(2)(343));                                                             
 
                tmr_registers(0)(345)    <= not(global_tmr_voter(0)(344));                                                             
                tmr_registers(1)(345)    <= not(global_tmr_voter(1)(344));                                                             
                tmr_registers(2)(345)    <= not(global_tmr_voter(2)(344));                                                             
 
                tmr_registers(0)(346)    <= not(global_tmr_voter(0)(345));                                                             
                tmr_registers(1)(346)    <= not(global_tmr_voter(1)(345));                                                             
                tmr_registers(2)(346)    <= not(global_tmr_voter(2)(345));                                                             
 
                tmr_registers(0)(347)    <= not(global_tmr_voter(0)(346));                                                             
                tmr_registers(1)(347)    <= not(global_tmr_voter(1)(346));                                                             
                tmr_registers(2)(347)    <= not(global_tmr_voter(2)(346));                                                             
 
                tmr_registers(0)(348)    <= not(global_tmr_voter(0)(347));                                                             
                tmr_registers(1)(348)    <= not(global_tmr_voter(1)(347));                                                             
                tmr_registers(2)(348)    <= not(global_tmr_voter(2)(347));                                                             
 
                tmr_registers(0)(349)    <= not(global_tmr_voter(0)(348));                                                             
                tmr_registers(1)(349)    <= not(global_tmr_voter(1)(348));                                                             
                tmr_registers(2)(349)    <= not(global_tmr_voter(2)(348));                                                             
 
                tmr_registers(0)(350)    <= not(global_tmr_voter(0)(349));                                                             
                tmr_registers(1)(350)    <= not(global_tmr_voter(1)(349));                                                             
                tmr_registers(2)(350)    <= not(global_tmr_voter(2)(349));                                                             
 
                tmr_registers(0)(351)    <= not(global_tmr_voter(0)(350));                                                             
                tmr_registers(1)(351)    <= not(global_tmr_voter(1)(350));                                                             
                tmr_registers(2)(351)    <= not(global_tmr_voter(2)(350));                                                             
 
                tmr_registers(0)(352)    <= not(global_tmr_voter(0)(351));                                                             
                tmr_registers(1)(352)    <= not(global_tmr_voter(1)(351));                                                             
                tmr_registers(2)(352)    <= not(global_tmr_voter(2)(351));                                                             
 
                tmr_registers(0)(353)    <= not(global_tmr_voter(0)(352));                                                             
                tmr_registers(1)(353)    <= not(global_tmr_voter(1)(352));                                                             
                tmr_registers(2)(353)    <= not(global_tmr_voter(2)(352));                                                             
 
                tmr_registers(0)(354)    <= not(global_tmr_voter(0)(353));                                                             
                tmr_registers(1)(354)    <= not(global_tmr_voter(1)(353));                                                             
                tmr_registers(2)(354)    <= not(global_tmr_voter(2)(353));                                                             
 
                tmr_registers(0)(355)    <= not(global_tmr_voter(0)(354));                                                             
                tmr_registers(1)(355)    <= not(global_tmr_voter(1)(354));                                                             
                tmr_registers(2)(355)    <= not(global_tmr_voter(2)(354));                                                             
 
                tmr_registers(0)(356)    <= not(global_tmr_voter(0)(355));                                                             
                tmr_registers(1)(356)    <= not(global_tmr_voter(1)(355));                                                             
                tmr_registers(2)(356)    <= not(global_tmr_voter(2)(355));                                                             
 
                tmr_registers(0)(357)    <= not(global_tmr_voter(0)(356));                                                             
                tmr_registers(1)(357)    <= not(global_tmr_voter(1)(356));                                                             
                tmr_registers(2)(357)    <= not(global_tmr_voter(2)(356));                                                             
 
                tmr_registers(0)(358)    <= not(global_tmr_voter(0)(357));                                                             
                tmr_registers(1)(358)    <= not(global_tmr_voter(1)(357));                                                             
                tmr_registers(2)(358)    <= not(global_tmr_voter(2)(357));                                                             
 
                tmr_registers(0)(359)    <= not(global_tmr_voter(0)(358));                                                             
                tmr_registers(1)(359)    <= not(global_tmr_voter(1)(358));                                                             
                tmr_registers(2)(359)    <= not(global_tmr_voter(2)(358));                                                             
 
                tmr_registers(0)(360)    <= not(global_tmr_voter(0)(359));                                                             
                tmr_registers(1)(360)    <= not(global_tmr_voter(1)(359));                                                             
                tmr_registers(2)(360)    <= not(global_tmr_voter(2)(359));                                                             
 
                tmr_registers(0)(361)    <= not(global_tmr_voter(0)(360));                                                             
                tmr_registers(1)(361)    <= not(global_tmr_voter(1)(360));                                                             
                tmr_registers(2)(361)    <= not(global_tmr_voter(2)(360));                                                             
 
                tmr_registers(0)(362)    <= not(global_tmr_voter(0)(361));                                                             
                tmr_registers(1)(362)    <= not(global_tmr_voter(1)(361));                                                             
                tmr_registers(2)(362)    <= not(global_tmr_voter(2)(361));                                                             
 
                tmr_registers(0)(363)    <= not(global_tmr_voter(0)(362));                                                             
                tmr_registers(1)(363)    <= not(global_tmr_voter(1)(362));                                                             
                tmr_registers(2)(363)    <= not(global_tmr_voter(2)(362));                                                             
 
                tmr_registers(0)(364)    <= not(global_tmr_voter(0)(363));                                                             
                tmr_registers(1)(364)    <= not(global_tmr_voter(1)(363));                                                             
                tmr_registers(2)(364)    <= not(global_tmr_voter(2)(363));                                                             
 
                tmr_registers(0)(365)    <= not(global_tmr_voter(0)(364));                                                             
                tmr_registers(1)(365)    <= not(global_tmr_voter(1)(364));                                                             
                tmr_registers(2)(365)    <= not(global_tmr_voter(2)(364));                                                             
 
                tmr_registers(0)(366)    <= not(global_tmr_voter(0)(365));                                                             
                tmr_registers(1)(366)    <= not(global_tmr_voter(1)(365));                                                             
                tmr_registers(2)(366)    <= not(global_tmr_voter(2)(365));                                                             
 
                tmr_registers(0)(367)    <= not(global_tmr_voter(0)(366));                                                             
                tmr_registers(1)(367)    <= not(global_tmr_voter(1)(366));                                                             
                tmr_registers(2)(367)    <= not(global_tmr_voter(2)(366));                                                             
 
                tmr_registers(0)(368)    <= not(global_tmr_voter(0)(367));                                                             
                tmr_registers(1)(368)    <= not(global_tmr_voter(1)(367));                                                             
                tmr_registers(2)(368)    <= not(global_tmr_voter(2)(367));                                                             
 
                tmr_registers(0)(369)    <= not(global_tmr_voter(0)(368));                                                             
                tmr_registers(1)(369)    <= not(global_tmr_voter(1)(368));                                                             
                tmr_registers(2)(369)    <= not(global_tmr_voter(2)(368));                                                             
 
                tmr_registers(0)(370)    <= not(global_tmr_voter(0)(369));                                                             
                tmr_registers(1)(370)    <= not(global_tmr_voter(1)(369));                                                             
                tmr_registers(2)(370)    <= not(global_tmr_voter(2)(369));                                                             
 
                tmr_registers(0)(371)    <= not(global_tmr_voter(0)(370));                                                             
                tmr_registers(1)(371)    <= not(global_tmr_voter(1)(370));                                                             
                tmr_registers(2)(371)    <= not(global_tmr_voter(2)(370));                                                             
 
                tmr_registers(0)(372)    <= not(global_tmr_voter(0)(371));                                                             
                tmr_registers(1)(372)    <= not(global_tmr_voter(1)(371));                                                             
                tmr_registers(2)(372)    <= not(global_tmr_voter(2)(371));                                                             
 
                tmr_registers(0)(373)    <= not(global_tmr_voter(0)(372));                                                             
                tmr_registers(1)(373)    <= not(global_tmr_voter(1)(372));                                                             
                tmr_registers(2)(373)    <= not(global_tmr_voter(2)(372));                                                             
 
                tmr_registers(0)(374)    <= not(global_tmr_voter(0)(373));                                                             
                tmr_registers(1)(374)    <= not(global_tmr_voter(1)(373));                                                             
                tmr_registers(2)(374)    <= not(global_tmr_voter(2)(373));                                                             
 
                tmr_registers(0)(375)    <= not(global_tmr_voter(0)(374));                                                             
                tmr_registers(1)(375)    <= not(global_tmr_voter(1)(374));                                                             
                tmr_registers(2)(375)    <= not(global_tmr_voter(2)(374));                                                             
 
                tmr_registers(0)(376)    <= not(global_tmr_voter(0)(375));                                                             
                tmr_registers(1)(376)    <= not(global_tmr_voter(1)(375));                                                             
                tmr_registers(2)(376)    <= not(global_tmr_voter(2)(375));                                                             
 
                tmr_registers(0)(377)    <= not(global_tmr_voter(0)(376));                                                             
                tmr_registers(1)(377)    <= not(global_tmr_voter(1)(376));                                                             
                tmr_registers(2)(377)    <= not(global_tmr_voter(2)(376));                                                             
 
                tmr_registers(0)(378)    <= not(global_tmr_voter(0)(377));                                                             
                tmr_registers(1)(378)    <= not(global_tmr_voter(1)(377));                                                             
                tmr_registers(2)(378)    <= not(global_tmr_voter(2)(377));                                                             
 
                tmr_registers(0)(379)    <= not(global_tmr_voter(0)(378));                                                             
                tmr_registers(1)(379)    <= not(global_tmr_voter(1)(378));                                                             
                tmr_registers(2)(379)    <= not(global_tmr_voter(2)(378));                                                             
 
                tmr_registers(0)(380)    <= not(global_tmr_voter(0)(379));                                                             
                tmr_registers(1)(380)    <= not(global_tmr_voter(1)(379));                                                             
                tmr_registers(2)(380)    <= not(global_tmr_voter(2)(379));                                                             
 
                tmr_registers(0)(381)    <= not(global_tmr_voter(0)(380));                                                             
                tmr_registers(1)(381)    <= not(global_tmr_voter(1)(380));                                                             
                tmr_registers(2)(381)    <= not(global_tmr_voter(2)(380));                                                             
 
                tmr_registers(0)(382)    <= not(global_tmr_voter(0)(381));                                                             
                tmr_registers(1)(382)    <= not(global_tmr_voter(1)(381));                                                             
                tmr_registers(2)(382)    <= not(global_tmr_voter(2)(381));                                                             
 
                tmr_registers(0)(383)    <= not(global_tmr_voter(0)(382));                                                             
                tmr_registers(1)(383)    <= not(global_tmr_voter(1)(382));                                                             
                tmr_registers(2)(383)    <= not(global_tmr_voter(2)(382));                                                             
 
                tmr_registers(0)(384)    <= not(global_tmr_voter(0)(383));                                                             
                tmr_registers(1)(384)    <= not(global_tmr_voter(1)(383));                                                             
                tmr_registers(2)(384)    <= not(global_tmr_voter(2)(383));                                                             
 
                tmr_registers(0)(385)    <= not(global_tmr_voter(0)(384));                                                             
                tmr_registers(1)(385)    <= not(global_tmr_voter(1)(384));                                                             
                tmr_registers(2)(385)    <= not(global_tmr_voter(2)(384));                                                             
 
                tmr_registers(0)(386)    <= not(global_tmr_voter(0)(385));                                                             
                tmr_registers(1)(386)    <= not(global_tmr_voter(1)(385));                                                             
                tmr_registers(2)(386)    <= not(global_tmr_voter(2)(385));                                                             
 
                tmr_registers(0)(387)    <= not(global_tmr_voter(0)(386));                                                             
                tmr_registers(1)(387)    <= not(global_tmr_voter(1)(386));                                                             
                tmr_registers(2)(387)    <= not(global_tmr_voter(2)(386));                                                             
 
                tmr_registers(0)(388)    <= not(global_tmr_voter(0)(387));                                                             
                tmr_registers(1)(388)    <= not(global_tmr_voter(1)(387));                                                             
                tmr_registers(2)(388)    <= not(global_tmr_voter(2)(387));                                                             
 
                tmr_registers(0)(389)    <= not(global_tmr_voter(0)(388));                                                             
                tmr_registers(1)(389)    <= not(global_tmr_voter(1)(388));                                                             
                tmr_registers(2)(389)    <= not(global_tmr_voter(2)(388));                                                             
 
                tmr_registers(0)(390)    <= not(global_tmr_voter(0)(389));                                                             
                tmr_registers(1)(390)    <= not(global_tmr_voter(1)(389));                                                             
                tmr_registers(2)(390)    <= not(global_tmr_voter(2)(389));                                                             
 
                tmr_registers(0)(391)    <= not(global_tmr_voter(0)(390));                                                             
                tmr_registers(1)(391)    <= not(global_tmr_voter(1)(390));                                                             
                tmr_registers(2)(391)    <= not(global_tmr_voter(2)(390));                                                             
 
                tmr_registers(0)(392)    <= not(global_tmr_voter(0)(391));                                                             
                tmr_registers(1)(392)    <= not(global_tmr_voter(1)(391));                                                             
                tmr_registers(2)(392)    <= not(global_tmr_voter(2)(391));                                                             
 
                tmr_registers(0)(393)    <= not(global_tmr_voter(0)(392));                                                             
                tmr_registers(1)(393)    <= not(global_tmr_voter(1)(392));                                                             
                tmr_registers(2)(393)    <= not(global_tmr_voter(2)(392));                                                             
 
                tmr_registers(0)(394)    <= not(global_tmr_voter(0)(393));                                                             
                tmr_registers(1)(394)    <= not(global_tmr_voter(1)(393));                                                             
                tmr_registers(2)(394)    <= not(global_tmr_voter(2)(393));                                                             
 
                tmr_registers(0)(395)    <= not(global_tmr_voter(0)(394));                                                             
                tmr_registers(1)(395)    <= not(global_tmr_voter(1)(394));                                                             
                tmr_registers(2)(395)    <= not(global_tmr_voter(2)(394));                                                             
 
                tmr_registers(0)(396)    <= not(global_tmr_voter(0)(395));                                                             
                tmr_registers(1)(396)    <= not(global_tmr_voter(1)(395));                                                             
                tmr_registers(2)(396)    <= not(global_tmr_voter(2)(395));                                                             
 
                tmr_registers(0)(397)    <= not(global_tmr_voter(0)(396));                                                             
                tmr_registers(1)(397)    <= not(global_tmr_voter(1)(396));                                                             
                tmr_registers(2)(397)    <= not(global_tmr_voter(2)(396));                                                             
 
                tmr_registers(0)(398)    <= not(global_tmr_voter(0)(397));                                                             
                tmr_registers(1)(398)    <= not(global_tmr_voter(1)(397));                                                             
                tmr_registers(2)(398)    <= not(global_tmr_voter(2)(397));                                                             
 
                tmr_registers(0)(399)    <= not(global_tmr_voter(0)(398));                                                             
                tmr_registers(1)(399)    <= not(global_tmr_voter(1)(398));                                                             
                tmr_registers(2)(399)    <= not(global_tmr_voter(2)(398));                                                             
 
                tmr_registers(0)(400)    <= not(global_tmr_voter(0)(399));                                                             
                tmr_registers(1)(400)    <= not(global_tmr_voter(1)(399));                                                             
                tmr_registers(2)(400)    <= not(global_tmr_voter(2)(399));                                                             
 
                tmr_registers(0)(401)    <= not(global_tmr_voter(0)(400));                                                             
                tmr_registers(1)(401)    <= not(global_tmr_voter(1)(400));                                                             
                tmr_registers(2)(401)    <= not(global_tmr_voter(2)(400));                                                             
 
                tmr_registers(0)(402)    <= not(global_tmr_voter(0)(401));                                                             
                tmr_registers(1)(402)    <= not(global_tmr_voter(1)(401));                                                             
                tmr_registers(2)(402)    <= not(global_tmr_voter(2)(401));                                                             
 
                tmr_registers(0)(403)    <= not(global_tmr_voter(0)(402));                                                             
                tmr_registers(1)(403)    <= not(global_tmr_voter(1)(402));                                                             
                tmr_registers(2)(403)    <= not(global_tmr_voter(2)(402));                                                             
 
                tmr_registers(0)(404)    <= not(global_tmr_voter(0)(403));                                                             
                tmr_registers(1)(404)    <= not(global_tmr_voter(1)(403));                                                             
                tmr_registers(2)(404)    <= not(global_tmr_voter(2)(403));                                                             
 
                tmr_registers(0)(405)    <= not(global_tmr_voter(0)(404));                                                             
                tmr_registers(1)(405)    <= not(global_tmr_voter(1)(404));                                                             
                tmr_registers(2)(405)    <= not(global_tmr_voter(2)(404));                                                             
 
                tmr_registers(0)(406)    <= not(global_tmr_voter(0)(405));                                                             
                tmr_registers(1)(406)    <= not(global_tmr_voter(1)(405));                                                             
                tmr_registers(2)(406)    <= not(global_tmr_voter(2)(405));                                                             
 
                tmr_registers(0)(407)    <= not(global_tmr_voter(0)(406));                                                             
                tmr_registers(1)(407)    <= not(global_tmr_voter(1)(406));                                                             
                tmr_registers(2)(407)    <= not(global_tmr_voter(2)(406));                                                             
 
                tmr_registers(0)(408)    <= not(global_tmr_voter(0)(407));                                                             
                tmr_registers(1)(408)    <= not(global_tmr_voter(1)(407));                                                             
                tmr_registers(2)(408)    <= not(global_tmr_voter(2)(407));                                                             
 
                tmr_registers(0)(409)    <= not(global_tmr_voter(0)(408));                                                             
                tmr_registers(1)(409)    <= not(global_tmr_voter(1)(408));                                                             
                tmr_registers(2)(409)    <= not(global_tmr_voter(2)(408));                                                             
 
                tmr_registers(0)(410)    <= not(global_tmr_voter(0)(409));                                                             
                tmr_registers(1)(410)    <= not(global_tmr_voter(1)(409));                                                             
                tmr_registers(2)(410)    <= not(global_tmr_voter(2)(409));                                                             
 
                tmr_registers(0)(411)    <= not(global_tmr_voter(0)(410));                                                             
                tmr_registers(1)(411)    <= not(global_tmr_voter(1)(410));                                                             
                tmr_registers(2)(411)    <= not(global_tmr_voter(2)(410));                                                             
 
                tmr_registers(0)(412)    <= not(global_tmr_voter(0)(411));                                                             
                tmr_registers(1)(412)    <= not(global_tmr_voter(1)(411));                                                             
                tmr_registers(2)(412)    <= not(global_tmr_voter(2)(411));                                                             
 
                tmr_registers(0)(413)    <= not(global_tmr_voter(0)(412));                                                             
                tmr_registers(1)(413)    <= not(global_tmr_voter(1)(412));                                                             
                tmr_registers(2)(413)    <= not(global_tmr_voter(2)(412));                                                             
 
                tmr_registers(0)(414)    <= not(global_tmr_voter(0)(413));                                                             
                tmr_registers(1)(414)    <= not(global_tmr_voter(1)(413));                                                             
                tmr_registers(2)(414)    <= not(global_tmr_voter(2)(413));                                                             
 
                tmr_registers(0)(415)    <= not(global_tmr_voter(0)(414));                                                             
                tmr_registers(1)(415)    <= not(global_tmr_voter(1)(414));                                                             
                tmr_registers(2)(415)    <= not(global_tmr_voter(2)(414));                                                             
 
                tmr_registers(0)(416)    <= not(global_tmr_voter(0)(415));                                                             
                tmr_registers(1)(416)    <= not(global_tmr_voter(1)(415));                                                             
                tmr_registers(2)(416)    <= not(global_tmr_voter(2)(415));                                                             
 
                tmr_registers(0)(417)    <= not(global_tmr_voter(0)(416));                                                             
                tmr_registers(1)(417)    <= not(global_tmr_voter(1)(416));                                                             
                tmr_registers(2)(417)    <= not(global_tmr_voter(2)(416));                                                             
 
                tmr_registers(0)(418)    <= not(global_tmr_voter(0)(417));                                                             
                tmr_registers(1)(418)    <= not(global_tmr_voter(1)(417));                                                             
                tmr_registers(2)(418)    <= not(global_tmr_voter(2)(417));                                                             
 
                tmr_registers(0)(419)    <= not(global_tmr_voter(0)(418));                                                             
                tmr_registers(1)(419)    <= not(global_tmr_voter(1)(418));                                                             
                tmr_registers(2)(419)    <= not(global_tmr_voter(2)(418));                                                             
 
                tmr_registers(0)(420)    <= not(global_tmr_voter(0)(419));                                                             
                tmr_registers(1)(420)    <= not(global_tmr_voter(1)(419));                                                             
                tmr_registers(2)(420)    <= not(global_tmr_voter(2)(419));                                                             
 
                tmr_registers(0)(421)    <= not(global_tmr_voter(0)(420));                                                             
                tmr_registers(1)(421)    <= not(global_tmr_voter(1)(420));                                                             
                tmr_registers(2)(421)    <= not(global_tmr_voter(2)(420));                                                             
 
                tmr_registers(0)(422)    <= not(global_tmr_voter(0)(421));                                                             
                tmr_registers(1)(422)    <= not(global_tmr_voter(1)(421));                                                             
                tmr_registers(2)(422)    <= not(global_tmr_voter(2)(421));                                                             
 
                tmr_registers(0)(423)    <= not(global_tmr_voter(0)(422));                                                             
                tmr_registers(1)(423)    <= not(global_tmr_voter(1)(422));                                                             
                tmr_registers(2)(423)    <= not(global_tmr_voter(2)(422));                                                             
 
                tmr_registers(0)(424)    <= not(global_tmr_voter(0)(423));                                                             
                tmr_registers(1)(424)    <= not(global_tmr_voter(1)(423));                                                             
                tmr_registers(2)(424)    <= not(global_tmr_voter(2)(423));                                                             
 
                tmr_registers(0)(425)    <= not(global_tmr_voter(0)(424));                                                             
                tmr_registers(1)(425)    <= not(global_tmr_voter(1)(424));                                                             
                tmr_registers(2)(425)    <= not(global_tmr_voter(2)(424));                                                             
 
                tmr_registers(0)(426)    <= not(global_tmr_voter(0)(425));                                                             
                tmr_registers(1)(426)    <= not(global_tmr_voter(1)(425));                                                             
                tmr_registers(2)(426)    <= not(global_tmr_voter(2)(425));                                                             
 
                tmr_registers(0)(427)    <= not(global_tmr_voter(0)(426));                                                             
                tmr_registers(1)(427)    <= not(global_tmr_voter(1)(426));                                                             
                tmr_registers(2)(427)    <= not(global_tmr_voter(2)(426));                                                             
 
                tmr_registers(0)(428)    <= not(global_tmr_voter(0)(427));                                                             
                tmr_registers(1)(428)    <= not(global_tmr_voter(1)(427));                                                             
                tmr_registers(2)(428)    <= not(global_tmr_voter(2)(427));                                                             
 
                tmr_registers(0)(429)    <= not(global_tmr_voter(0)(428));                                                             
                tmr_registers(1)(429)    <= not(global_tmr_voter(1)(428));                                                             
                tmr_registers(2)(429)    <= not(global_tmr_voter(2)(428));                                                             
 
                tmr_registers(0)(430)    <= not(global_tmr_voter(0)(429));                                                             
                tmr_registers(1)(430)    <= not(global_tmr_voter(1)(429));                                                             
                tmr_registers(2)(430)    <= not(global_tmr_voter(2)(429));                                                             
 
                tmr_registers(0)(431)    <= not(global_tmr_voter(0)(430));                                                             
                tmr_registers(1)(431)    <= not(global_tmr_voter(1)(430));                                                             
                tmr_registers(2)(431)    <= not(global_tmr_voter(2)(430));                                                             
 
                tmr_registers(0)(432)    <= not(global_tmr_voter(0)(431));                                                             
                tmr_registers(1)(432)    <= not(global_tmr_voter(1)(431));                                                             
                tmr_registers(2)(432)    <= not(global_tmr_voter(2)(431));                                                             
 
                tmr_registers(0)(433)    <= not(global_tmr_voter(0)(432));                                                             
                tmr_registers(1)(433)    <= not(global_tmr_voter(1)(432));                                                             
                tmr_registers(2)(433)    <= not(global_tmr_voter(2)(432));                                                             
 
                tmr_registers(0)(434)    <= not(global_tmr_voter(0)(433));                                                             
                tmr_registers(1)(434)    <= not(global_tmr_voter(1)(433));                                                             
                tmr_registers(2)(434)    <= not(global_tmr_voter(2)(433));                                                             
 
                tmr_registers(0)(435)    <= not(global_tmr_voter(0)(434));                                                             
                tmr_registers(1)(435)    <= not(global_tmr_voter(1)(434));                                                             
                tmr_registers(2)(435)    <= not(global_tmr_voter(2)(434));                                                             
 
                tmr_registers(0)(436)    <= not(global_tmr_voter(0)(435));                                                             
                tmr_registers(1)(436)    <= not(global_tmr_voter(1)(435));                                                             
                tmr_registers(2)(436)    <= not(global_tmr_voter(2)(435));                                                             
 
                tmr_registers(0)(437)    <= not(global_tmr_voter(0)(436));                                                             
                tmr_registers(1)(437)    <= not(global_tmr_voter(1)(436));                                                             
                tmr_registers(2)(437)    <= not(global_tmr_voter(2)(436));                                                             
 
                tmr_registers(0)(438)    <= not(global_tmr_voter(0)(437));                                                             
                tmr_registers(1)(438)    <= not(global_tmr_voter(1)(437));                                                             
                tmr_registers(2)(438)    <= not(global_tmr_voter(2)(437));                                                             
 
                tmr_registers(0)(439)    <= not(global_tmr_voter(0)(438));                                                             
                tmr_registers(1)(439)    <= not(global_tmr_voter(1)(438));                                                             
                tmr_registers(2)(439)    <= not(global_tmr_voter(2)(438));                                                             
 
                tmr_registers(0)(440)    <= not(global_tmr_voter(0)(439));                                                             
                tmr_registers(1)(440)    <= not(global_tmr_voter(1)(439));                                                             
                tmr_registers(2)(440)    <= not(global_tmr_voter(2)(439));                                                             
 
                tmr_registers(0)(441)    <= not(global_tmr_voter(0)(440));                                                             
                tmr_registers(1)(441)    <= not(global_tmr_voter(1)(440));                                                             
                tmr_registers(2)(441)    <= not(global_tmr_voter(2)(440));                                                             
 
                tmr_registers(0)(442)    <= not(global_tmr_voter(0)(441));                                                             
                tmr_registers(1)(442)    <= not(global_tmr_voter(1)(441));                                                             
                tmr_registers(2)(442)    <= not(global_tmr_voter(2)(441));                                                             
 
                tmr_registers(0)(443)    <= not(global_tmr_voter(0)(442));                                                             
                tmr_registers(1)(443)    <= not(global_tmr_voter(1)(442));                                                             
                tmr_registers(2)(443)    <= not(global_tmr_voter(2)(442));                                                             
 
                tmr_registers(0)(444)    <= not(global_tmr_voter(0)(443));                                                             
                tmr_registers(1)(444)    <= not(global_tmr_voter(1)(443));                                                             
                tmr_registers(2)(444)    <= not(global_tmr_voter(2)(443));                                                             
 
                tmr_registers(0)(445)    <= not(global_tmr_voter(0)(444));                                                             
                tmr_registers(1)(445)    <= not(global_tmr_voter(1)(444));                                                             
                tmr_registers(2)(445)    <= not(global_tmr_voter(2)(444));                                                             
 
                tmr_registers(0)(446)    <= not(global_tmr_voter(0)(445));                                                             
                tmr_registers(1)(446)    <= not(global_tmr_voter(1)(445));                                                             
                tmr_registers(2)(446)    <= not(global_tmr_voter(2)(445));                                                             
 
                tmr_registers(0)(447)    <= not(global_tmr_voter(0)(446));                                                             
                tmr_registers(1)(447)    <= not(global_tmr_voter(1)(446));                                                             
                tmr_registers(2)(447)    <= not(global_tmr_voter(2)(446));                                                             
 
                tmr_registers(0)(448)    <= not(global_tmr_voter(0)(447));                                                             
                tmr_registers(1)(448)    <= not(global_tmr_voter(1)(447));                                                             
                tmr_registers(2)(448)    <= not(global_tmr_voter(2)(447));                                                             
 
                tmr_registers(0)(449)    <= not(global_tmr_voter(0)(448));                                                             
                tmr_registers(1)(449)    <= not(global_tmr_voter(1)(448));                                                             
                tmr_registers(2)(449)    <= not(global_tmr_voter(2)(448));                                                             
 
                tmr_registers(0)(450)    <= not(global_tmr_voter(0)(449));                                                             
                tmr_registers(1)(450)    <= not(global_tmr_voter(1)(449));                                                             
                tmr_registers(2)(450)    <= not(global_tmr_voter(2)(449));                                                             
 
                tmr_registers(0)(451)    <= not(global_tmr_voter(0)(450));                                                             
                tmr_registers(1)(451)    <= not(global_tmr_voter(1)(450));                                                             
                tmr_registers(2)(451)    <= not(global_tmr_voter(2)(450));                                                             
 
                tmr_registers(0)(452)    <= not(global_tmr_voter(0)(451));                                                             
                tmr_registers(1)(452)    <= not(global_tmr_voter(1)(451));                                                             
                tmr_registers(2)(452)    <= not(global_tmr_voter(2)(451));                                                             
 
                tmr_registers(0)(453)    <= not(global_tmr_voter(0)(452));                                                             
                tmr_registers(1)(453)    <= not(global_tmr_voter(1)(452));                                                             
                tmr_registers(2)(453)    <= not(global_tmr_voter(2)(452));                                                             
 
                tmr_registers(0)(454)    <= not(global_tmr_voter(0)(453));                                                             
                tmr_registers(1)(454)    <= not(global_tmr_voter(1)(453));                                                             
                tmr_registers(2)(454)    <= not(global_tmr_voter(2)(453));                                                             
 
                tmr_registers(0)(455)    <= not(global_tmr_voter(0)(454));                                                             
                tmr_registers(1)(455)    <= not(global_tmr_voter(1)(454));                                                             
                tmr_registers(2)(455)    <= not(global_tmr_voter(2)(454));                                                             
 
                tmr_registers(0)(456)    <= not(global_tmr_voter(0)(455));                                                             
                tmr_registers(1)(456)    <= not(global_tmr_voter(1)(455));                                                             
                tmr_registers(2)(456)    <= not(global_tmr_voter(2)(455));                                                             
 
                tmr_registers(0)(457)    <= not(global_tmr_voter(0)(456));                                                             
                tmr_registers(1)(457)    <= not(global_tmr_voter(1)(456));                                                             
                tmr_registers(2)(457)    <= not(global_tmr_voter(2)(456));                                                             
 
                tmr_registers(0)(458)    <= not(global_tmr_voter(0)(457));                                                             
                tmr_registers(1)(458)    <= not(global_tmr_voter(1)(457));                                                             
                tmr_registers(2)(458)    <= not(global_tmr_voter(2)(457));                                                             
 
                tmr_registers(0)(459)    <= not(global_tmr_voter(0)(458));                                                             
                tmr_registers(1)(459)    <= not(global_tmr_voter(1)(458));                                                             
                tmr_registers(2)(459)    <= not(global_tmr_voter(2)(458));                                                             
 
                tmr_registers(0)(460)    <= not(global_tmr_voter(0)(459));                                                             
                tmr_registers(1)(460)    <= not(global_tmr_voter(1)(459));                                                             
                tmr_registers(2)(460)    <= not(global_tmr_voter(2)(459));                                                             
 
                tmr_registers(0)(461)    <= not(global_tmr_voter(0)(460));                                                             
                tmr_registers(1)(461)    <= not(global_tmr_voter(1)(460));                                                             
                tmr_registers(2)(461)    <= not(global_tmr_voter(2)(460));                                                             
 
                tmr_registers(0)(462)    <= not(global_tmr_voter(0)(461));                                                             
                tmr_registers(1)(462)    <= not(global_tmr_voter(1)(461));                                                             
                tmr_registers(2)(462)    <= not(global_tmr_voter(2)(461));                                                             
 
                tmr_registers(0)(463)    <= not(global_tmr_voter(0)(462));                                                             
                tmr_registers(1)(463)    <= not(global_tmr_voter(1)(462));                                                             
                tmr_registers(2)(463)    <= not(global_tmr_voter(2)(462));                                                             
 
                tmr_registers(0)(464)    <= not(global_tmr_voter(0)(463));                                                             
                tmr_registers(1)(464)    <= not(global_tmr_voter(1)(463));                                                             
                tmr_registers(2)(464)    <= not(global_tmr_voter(2)(463));                                                             
 
                tmr_registers(0)(465)    <= not(global_tmr_voter(0)(464));                                                             
                tmr_registers(1)(465)    <= not(global_tmr_voter(1)(464));                                                             
                tmr_registers(2)(465)    <= not(global_tmr_voter(2)(464));                                                             
 
                tmr_registers(0)(466)    <= not(global_tmr_voter(0)(465));                                                             
                tmr_registers(1)(466)    <= not(global_tmr_voter(1)(465));                                                             
                tmr_registers(2)(466)    <= not(global_tmr_voter(2)(465));                                                             
 
                tmr_registers(0)(467)    <= not(global_tmr_voter(0)(466));                                                             
                tmr_registers(1)(467)    <= not(global_tmr_voter(1)(466));                                                             
                tmr_registers(2)(467)    <= not(global_tmr_voter(2)(466));                                                             
 
                tmr_registers(0)(468)    <= not(global_tmr_voter(0)(467));                                                             
                tmr_registers(1)(468)    <= not(global_tmr_voter(1)(467));                                                             
                tmr_registers(2)(468)    <= not(global_tmr_voter(2)(467));                                                             
 
                tmr_registers(0)(469)    <= not(global_tmr_voter(0)(468));                                                             
                tmr_registers(1)(469)    <= not(global_tmr_voter(1)(468));                                                             
                tmr_registers(2)(469)    <= not(global_tmr_voter(2)(468));                                                             
 
                tmr_registers(0)(470)    <= not(global_tmr_voter(0)(469));                                                             
                tmr_registers(1)(470)    <= not(global_tmr_voter(1)(469));                                                             
                tmr_registers(2)(470)    <= not(global_tmr_voter(2)(469));                                                             
 
                tmr_registers(0)(471)    <= not(global_tmr_voter(0)(470));                                                             
                tmr_registers(1)(471)    <= not(global_tmr_voter(1)(470));                                                             
                tmr_registers(2)(471)    <= not(global_tmr_voter(2)(470));                                                             
 
                tmr_registers(0)(472)    <= not(global_tmr_voter(0)(471));                                                             
                tmr_registers(1)(472)    <= not(global_tmr_voter(1)(471));                                                             
                tmr_registers(2)(472)    <= not(global_tmr_voter(2)(471));                                                             
 
                tmr_registers(0)(473)    <= not(global_tmr_voter(0)(472));                                                             
                tmr_registers(1)(473)    <= not(global_tmr_voter(1)(472));                                                             
                tmr_registers(2)(473)    <= not(global_tmr_voter(2)(472));                                                             
 
                tmr_registers(0)(474)    <= not(global_tmr_voter(0)(473));                                                             
                tmr_registers(1)(474)    <= not(global_tmr_voter(1)(473));                                                             
                tmr_registers(2)(474)    <= not(global_tmr_voter(2)(473));                                                             
 
                tmr_registers(0)(475)    <= not(global_tmr_voter(0)(474));                                                             
                tmr_registers(1)(475)    <= not(global_tmr_voter(1)(474));                                                             
                tmr_registers(2)(475)    <= not(global_tmr_voter(2)(474));                                                             
 
                tmr_registers(0)(476)    <= not(global_tmr_voter(0)(475));                                                             
                tmr_registers(1)(476)    <= not(global_tmr_voter(1)(475));                                                             
                tmr_registers(2)(476)    <= not(global_tmr_voter(2)(475));                                                             
 
                tmr_registers(0)(477)    <= not(global_tmr_voter(0)(476));                                                             
                tmr_registers(1)(477)    <= not(global_tmr_voter(1)(476));                                                             
                tmr_registers(2)(477)    <= not(global_tmr_voter(2)(476));                                                             
 
                tmr_registers(0)(478)    <= not(global_tmr_voter(0)(477));                                                             
                tmr_registers(1)(478)    <= not(global_tmr_voter(1)(477));                                                             
                tmr_registers(2)(478)    <= not(global_tmr_voter(2)(477));                                                             
 
                tmr_registers(0)(479)    <= not(global_tmr_voter(0)(478));                                                             
                tmr_registers(1)(479)    <= not(global_tmr_voter(1)(478));                                                             
                tmr_registers(2)(479)    <= not(global_tmr_voter(2)(478));                                                             
 
                tmr_registers(0)(480)    <= not(global_tmr_voter(0)(479));                                                             
                tmr_registers(1)(480)    <= not(global_tmr_voter(1)(479));                                                             
                tmr_registers(2)(480)    <= not(global_tmr_voter(2)(479));                                                             
 
                tmr_registers(0)(481)    <= not(global_tmr_voter(0)(480));                                                             
                tmr_registers(1)(481)    <= not(global_tmr_voter(1)(480));                                                             
                tmr_registers(2)(481)    <= not(global_tmr_voter(2)(480));                                                             
 
                tmr_registers(0)(482)    <= not(global_tmr_voter(0)(481));                                                             
                tmr_registers(1)(482)    <= not(global_tmr_voter(1)(481));                                                             
                tmr_registers(2)(482)    <= not(global_tmr_voter(2)(481));                                                             
 
                tmr_registers(0)(483)    <= not(global_tmr_voter(0)(482));                                                             
                tmr_registers(1)(483)    <= not(global_tmr_voter(1)(482));                                                             
                tmr_registers(2)(483)    <= not(global_tmr_voter(2)(482));                                                             
 
                tmr_registers(0)(484)    <= not(global_tmr_voter(0)(483));                                                             
                tmr_registers(1)(484)    <= not(global_tmr_voter(1)(483));                                                             
                tmr_registers(2)(484)    <= not(global_tmr_voter(2)(483));                                                             
 
                tmr_registers(0)(485)    <= not(global_tmr_voter(0)(484));                                                             
                tmr_registers(1)(485)    <= not(global_tmr_voter(1)(484));                                                             
                tmr_registers(2)(485)    <= not(global_tmr_voter(2)(484));                                                             
 
                tmr_registers(0)(486)    <= not(global_tmr_voter(0)(485));                                                             
                tmr_registers(1)(486)    <= not(global_tmr_voter(1)(485));                                                             
                tmr_registers(2)(486)    <= not(global_tmr_voter(2)(485));                                                             
 
                tmr_registers(0)(487)    <= not(global_tmr_voter(0)(486));                                                             
                tmr_registers(1)(487)    <= not(global_tmr_voter(1)(486));                                                             
                tmr_registers(2)(487)    <= not(global_tmr_voter(2)(486));                                                             
 
                tmr_registers(0)(488)    <= not(global_tmr_voter(0)(487));                                                             
                tmr_registers(1)(488)    <= not(global_tmr_voter(1)(487));                                                             
                tmr_registers(2)(488)    <= not(global_tmr_voter(2)(487));                                                             
 
                tmr_registers(0)(489)    <= not(global_tmr_voter(0)(488));                                                             
                tmr_registers(1)(489)    <= not(global_tmr_voter(1)(488));                                                             
                tmr_registers(2)(489)    <= not(global_tmr_voter(2)(488));                                                             
 
                tmr_registers(0)(490)    <= not(global_tmr_voter(0)(489));                                                             
                tmr_registers(1)(490)    <= not(global_tmr_voter(1)(489));                                                             
                tmr_registers(2)(490)    <= not(global_tmr_voter(2)(489));                                                             
 
                tmr_registers(0)(491)    <= not(global_tmr_voter(0)(490));                                                             
                tmr_registers(1)(491)    <= not(global_tmr_voter(1)(490));                                                             
                tmr_registers(2)(491)    <= not(global_tmr_voter(2)(490));                                                             
 
                tmr_registers(0)(492)    <= not(global_tmr_voter(0)(491));                                                             
                tmr_registers(1)(492)    <= not(global_tmr_voter(1)(491));                                                             
                tmr_registers(2)(492)    <= not(global_tmr_voter(2)(491));                                                             
 
                tmr_registers(0)(493)    <= not(global_tmr_voter(0)(492));                                                             
                tmr_registers(1)(493)    <= not(global_tmr_voter(1)(492));                                                             
                tmr_registers(2)(493)    <= not(global_tmr_voter(2)(492));                                                             
 
                tmr_registers(0)(494)    <= not(global_tmr_voter(0)(493));                                                             
                tmr_registers(1)(494)    <= not(global_tmr_voter(1)(493));                                                             
                tmr_registers(2)(494)    <= not(global_tmr_voter(2)(493));                                                             
 
                tmr_registers(0)(495)    <= not(global_tmr_voter(0)(494));                                                             
                tmr_registers(1)(495)    <= not(global_tmr_voter(1)(494));                                                             
                tmr_registers(2)(495)    <= not(global_tmr_voter(2)(494));                                                             
 
                tmr_registers(0)(496)    <= not(global_tmr_voter(0)(495));                                                             
                tmr_registers(1)(496)    <= not(global_tmr_voter(1)(495));                                                             
                tmr_registers(2)(496)    <= not(global_tmr_voter(2)(495));                                                             
 
                tmr_registers(0)(497)    <= not(global_tmr_voter(0)(496));                                                             
                tmr_registers(1)(497)    <= not(global_tmr_voter(1)(496));                                                             
                tmr_registers(2)(497)    <= not(global_tmr_voter(2)(496));                                                             
 
                tmr_registers(0)(498)    <= not(global_tmr_voter(0)(497));                                                             
                tmr_registers(1)(498)    <= not(global_tmr_voter(1)(497));                                                             
                tmr_registers(2)(498)    <= not(global_tmr_voter(2)(497));                                                             
 
                tmr_registers(0)(499)    <= not(global_tmr_voter(0)(498));                                                             
                tmr_registers(1)(499)    <= not(global_tmr_voter(1)(498));                                                             
                tmr_registers(2)(499)    <= not(global_tmr_voter(2)(498));                                                             
 
                tmr_registers(0)(500)    <= not(global_tmr_voter(0)(499));                                                             
                tmr_registers(1)(500)    <= not(global_tmr_voter(1)(499));                                                             
                tmr_registers(2)(500)    <= not(global_tmr_voter(2)(499));                                                             
 
                tmr_registers(0)(501)    <= not(global_tmr_voter(0)(500));                                                             
                tmr_registers(1)(501)    <= not(global_tmr_voter(1)(500));                                                             
                tmr_registers(2)(501)    <= not(global_tmr_voter(2)(500));                                                             
 
                tmr_registers(0)(502)    <= not(global_tmr_voter(0)(501));                                                             
                tmr_registers(1)(502)    <= not(global_tmr_voter(1)(501));                                                             
                tmr_registers(2)(502)    <= not(global_tmr_voter(2)(501));                                                             
 
                tmr_registers(0)(503)    <= not(global_tmr_voter(0)(502));                                                             
                tmr_registers(1)(503)    <= not(global_tmr_voter(1)(502));                                                             
                tmr_registers(2)(503)    <= not(global_tmr_voter(2)(502));                                                             
 
                tmr_registers(0)(504)    <= not(global_tmr_voter(0)(503));                                                             
                tmr_registers(1)(504)    <= not(global_tmr_voter(1)(503));                                                             
                tmr_registers(2)(504)    <= not(global_tmr_voter(2)(503));                                                             
 
                tmr_registers(0)(505)    <= not(global_tmr_voter(0)(504));                                                             
                tmr_registers(1)(505)    <= not(global_tmr_voter(1)(504));                                                             
                tmr_registers(2)(505)    <= not(global_tmr_voter(2)(504));                                                             
 
                tmr_registers(0)(506)    <= not(global_tmr_voter(0)(505));                                                             
                tmr_registers(1)(506)    <= not(global_tmr_voter(1)(505));                                                             
                tmr_registers(2)(506)    <= not(global_tmr_voter(2)(505));                                                             
 
                tmr_registers(0)(507)    <= not(global_tmr_voter(0)(506));                                                             
                tmr_registers(1)(507)    <= not(global_tmr_voter(1)(506));                                                             
                tmr_registers(2)(507)    <= not(global_tmr_voter(2)(506));                                                             
 
                tmr_registers(0)(508)    <= not(global_tmr_voter(0)(507));                                                             
                tmr_registers(1)(508)    <= not(global_tmr_voter(1)(507));                                                             
                tmr_registers(2)(508)    <= not(global_tmr_voter(2)(507));                                                             
 
                tmr_registers(0)(509)    <= not(global_tmr_voter(0)(508));                                                             
                tmr_registers(1)(509)    <= not(global_tmr_voter(1)(508));                                                             
                tmr_registers(2)(509)    <= not(global_tmr_voter(2)(508));                                                             
 
                tmr_registers(0)(510)    <= not(global_tmr_voter(0)(509));                                                             
                tmr_registers(1)(510)    <= not(global_tmr_voter(1)(509));                                                             
                tmr_registers(2)(510)    <= not(global_tmr_voter(2)(509));                                                             
 
                tmr_registers(0)(511)    <= not(global_tmr_voter(0)(510));                                                             
                tmr_registers(1)(511)    <= not(global_tmr_voter(1)(510));                                                             
                tmr_registers(2)(511)    <= not(global_tmr_voter(2)(510));                                                             
 
                tmr_registers(0)(512)    <= not(global_tmr_voter(0)(511));                                                             
                tmr_registers(1)(512)    <= not(global_tmr_voter(1)(511));                                                             
                tmr_registers(2)(512)    <= not(global_tmr_voter(2)(511));                                                             
 
                tmr_registers(0)(513)    <= not(global_tmr_voter(0)(512));                                                             
                tmr_registers(1)(513)    <= not(global_tmr_voter(1)(512));                                                             
                tmr_registers(2)(513)    <= not(global_tmr_voter(2)(512));                                                             
 
                tmr_registers(0)(514)    <= not(global_tmr_voter(0)(513));                                                             
                tmr_registers(1)(514)    <= not(global_tmr_voter(1)(513));                                                             
                tmr_registers(2)(514)    <= not(global_tmr_voter(2)(513));                                                             
 
                tmr_registers(0)(515)    <= not(global_tmr_voter(0)(514));                                                             
                tmr_registers(1)(515)    <= not(global_tmr_voter(1)(514));                                                             
                tmr_registers(2)(515)    <= not(global_tmr_voter(2)(514));                                                             
 
                tmr_registers(0)(516)    <= not(global_tmr_voter(0)(515));                                                             
                tmr_registers(1)(516)    <= not(global_tmr_voter(1)(515));                                                             
                tmr_registers(2)(516)    <= not(global_tmr_voter(2)(515));                                                             
 
                tmr_registers(0)(517)    <= not(global_tmr_voter(0)(516));                                                             
                tmr_registers(1)(517)    <= not(global_tmr_voter(1)(516));                                                             
                tmr_registers(2)(517)    <= not(global_tmr_voter(2)(516));                                                             
 
                tmr_registers(0)(518)    <= not(global_tmr_voter(0)(517));                                                             
                tmr_registers(1)(518)    <= not(global_tmr_voter(1)(517));                                                             
                tmr_registers(2)(518)    <= not(global_tmr_voter(2)(517));                                                             
 
                tmr_registers(0)(519)    <= not(global_tmr_voter(0)(518));                                                             
                tmr_registers(1)(519)    <= not(global_tmr_voter(1)(518));                                                             
                tmr_registers(2)(519)    <= not(global_tmr_voter(2)(518));                                                             
 
                tmr_registers(0)(520)    <= not(global_tmr_voter(0)(519));                                                             
                tmr_registers(1)(520)    <= not(global_tmr_voter(1)(519));                                                             
                tmr_registers(2)(520)    <= not(global_tmr_voter(2)(519));                                                             
 
                tmr_registers(0)(521)    <= not(global_tmr_voter(0)(520));                                                             
                tmr_registers(1)(521)    <= not(global_tmr_voter(1)(520));                                                             
                tmr_registers(2)(521)    <= not(global_tmr_voter(2)(520));                                                             
 
                tmr_registers(0)(522)    <= not(global_tmr_voter(0)(521));                                                             
                tmr_registers(1)(522)    <= not(global_tmr_voter(1)(521));                                                             
                tmr_registers(2)(522)    <= not(global_tmr_voter(2)(521));                                                             
 
                tmr_registers(0)(523)    <= not(global_tmr_voter(0)(522));                                                             
                tmr_registers(1)(523)    <= not(global_tmr_voter(1)(522));                                                             
                tmr_registers(2)(523)    <= not(global_tmr_voter(2)(522));                                                             
 
                tmr_registers(0)(524)    <= not(global_tmr_voter(0)(523));                                                             
                tmr_registers(1)(524)    <= not(global_tmr_voter(1)(523));                                                             
                tmr_registers(2)(524)    <= not(global_tmr_voter(2)(523));                                                             
 
                tmr_registers(0)(525)    <= not(global_tmr_voter(0)(524));                                                             
                tmr_registers(1)(525)    <= not(global_tmr_voter(1)(524));                                                             
                tmr_registers(2)(525)    <= not(global_tmr_voter(2)(524));                                                             
 
                tmr_registers(0)(526)    <= not(global_tmr_voter(0)(525));                                                             
                tmr_registers(1)(526)    <= not(global_tmr_voter(1)(525));                                                             
                tmr_registers(2)(526)    <= not(global_tmr_voter(2)(525));                                                             
 
                tmr_registers(0)(527)    <= not(global_tmr_voter(0)(526));                                                             
                tmr_registers(1)(527)    <= not(global_tmr_voter(1)(526));                                                             
                tmr_registers(2)(527)    <= not(global_tmr_voter(2)(526));                                                             
 
                tmr_registers(0)(528)    <= not(global_tmr_voter(0)(527));                                                             
                tmr_registers(1)(528)    <= not(global_tmr_voter(1)(527));                                                             
                tmr_registers(2)(528)    <= not(global_tmr_voter(2)(527));                                                             
 
                tmr_registers(0)(529)    <= not(global_tmr_voter(0)(528));                                                             
                tmr_registers(1)(529)    <= not(global_tmr_voter(1)(528));                                                             
                tmr_registers(2)(529)    <= not(global_tmr_voter(2)(528));                                                             
 
                tmr_registers(0)(530)    <= not(global_tmr_voter(0)(529));                                                             
                tmr_registers(1)(530)    <= not(global_tmr_voter(1)(529));                                                             
                tmr_registers(2)(530)    <= not(global_tmr_voter(2)(529));                                                             
 
                tmr_registers(0)(531)    <= not(global_tmr_voter(0)(530));                                                             
                tmr_registers(1)(531)    <= not(global_tmr_voter(1)(530));                                                             
                tmr_registers(2)(531)    <= not(global_tmr_voter(2)(530));                                                             
 
                tmr_registers(0)(532)    <= not(global_tmr_voter(0)(531));                                                             
                tmr_registers(1)(532)    <= not(global_tmr_voter(1)(531));                                                             
                tmr_registers(2)(532)    <= not(global_tmr_voter(2)(531));                                                             
 
                tmr_registers(0)(533)    <= not(global_tmr_voter(0)(532));                                                             
                tmr_registers(1)(533)    <= not(global_tmr_voter(1)(532));                                                             
                tmr_registers(2)(533)    <= not(global_tmr_voter(2)(532));                                                             
 
                tmr_registers(0)(534)    <= not(global_tmr_voter(0)(533));                                                             
                tmr_registers(1)(534)    <= not(global_tmr_voter(1)(533));                                                             
                tmr_registers(2)(534)    <= not(global_tmr_voter(2)(533));                                                             
 
                tmr_registers(0)(535)    <= not(global_tmr_voter(0)(534));                                                             
                tmr_registers(1)(535)    <= not(global_tmr_voter(1)(534));                                                             
                tmr_registers(2)(535)    <= not(global_tmr_voter(2)(534));                                                             
 
                tmr_registers(0)(536)    <= not(global_tmr_voter(0)(535));                                                             
                tmr_registers(1)(536)    <= not(global_tmr_voter(1)(535));                                                             
                tmr_registers(2)(536)    <= not(global_tmr_voter(2)(535));                                                             
 
                tmr_registers(0)(537)    <= not(global_tmr_voter(0)(536));                                                             
                tmr_registers(1)(537)    <= not(global_tmr_voter(1)(536));                                                             
                tmr_registers(2)(537)    <= not(global_tmr_voter(2)(536));                                                             
 
                tmr_registers(0)(538)    <= not(global_tmr_voter(0)(537));                                                             
                tmr_registers(1)(538)    <= not(global_tmr_voter(1)(537));                                                             
                tmr_registers(2)(538)    <= not(global_tmr_voter(2)(537));                                                             
 
                tmr_registers(0)(539)    <= not(global_tmr_voter(0)(538));                                                             
                tmr_registers(1)(539)    <= not(global_tmr_voter(1)(538));                                                             
                tmr_registers(2)(539)    <= not(global_tmr_voter(2)(538));                                                             
 
                tmr_registers(0)(540)    <= not(global_tmr_voter(0)(539));                                                             
                tmr_registers(1)(540)    <= not(global_tmr_voter(1)(539));                                                             
                tmr_registers(2)(540)    <= not(global_tmr_voter(2)(539));                                                             
 
                tmr_registers(0)(541)    <= not(global_tmr_voter(0)(540));                                                             
                tmr_registers(1)(541)    <= not(global_tmr_voter(1)(540));                                                             
                tmr_registers(2)(541)    <= not(global_tmr_voter(2)(540));                                                             
 
                tmr_registers(0)(542)    <= not(global_tmr_voter(0)(541));                                                             
                tmr_registers(1)(542)    <= not(global_tmr_voter(1)(541));                                                             
                tmr_registers(2)(542)    <= not(global_tmr_voter(2)(541));                                                             
 
                tmr_registers(0)(543)    <= not(global_tmr_voter(0)(542));                                                             
                tmr_registers(1)(543)    <= not(global_tmr_voter(1)(542));                                                             
                tmr_registers(2)(543)    <= not(global_tmr_voter(2)(542));                                                             
 
                tmr_registers(0)(544)    <= not(global_tmr_voter(0)(543));                                                             
                tmr_registers(1)(544)    <= not(global_tmr_voter(1)(543));                                                             
                tmr_registers(2)(544)    <= not(global_tmr_voter(2)(543));                                                             
 
                tmr_registers(0)(545)    <= not(global_tmr_voter(0)(544));                                                             
                tmr_registers(1)(545)    <= not(global_tmr_voter(1)(544));                                                             
                tmr_registers(2)(545)    <= not(global_tmr_voter(2)(544));                                                             
 
                tmr_registers(0)(546)    <= not(global_tmr_voter(0)(545));                                                             
                tmr_registers(1)(546)    <= not(global_tmr_voter(1)(545));                                                             
                tmr_registers(2)(546)    <= not(global_tmr_voter(2)(545));                                                             
 
                tmr_registers(0)(547)    <= not(global_tmr_voter(0)(546));                                                             
                tmr_registers(1)(547)    <= not(global_tmr_voter(1)(546));                                                             
                tmr_registers(2)(547)    <= not(global_tmr_voter(2)(546));                                                             
 
                tmr_registers(0)(548)    <= not(global_tmr_voter(0)(547));                                                             
                tmr_registers(1)(548)    <= not(global_tmr_voter(1)(547));                                                             
                tmr_registers(2)(548)    <= not(global_tmr_voter(2)(547));                                                             
 
                tmr_registers(0)(549)    <= not(global_tmr_voter(0)(548));                                                             
                tmr_registers(1)(549)    <= not(global_tmr_voter(1)(548));                                                             
                tmr_registers(2)(549)    <= not(global_tmr_voter(2)(548));                                                             
 
                tmr_registers(0)(550)    <= not(global_tmr_voter(0)(549));                                                             
                tmr_registers(1)(550)    <= not(global_tmr_voter(1)(549));                                                             
                tmr_registers(2)(550)    <= not(global_tmr_voter(2)(549));                                                             
 
                tmr_registers(0)(551)    <= not(global_tmr_voter(0)(550));                                                             
                tmr_registers(1)(551)    <= not(global_tmr_voter(1)(550));                                                             
                tmr_registers(2)(551)    <= not(global_tmr_voter(2)(550));                                                             
 
                tmr_registers(0)(552)    <= not(global_tmr_voter(0)(551));                                                             
                tmr_registers(1)(552)    <= not(global_tmr_voter(1)(551));                                                             
                tmr_registers(2)(552)    <= not(global_tmr_voter(2)(551));                                                             
 
                tmr_registers(0)(553)    <= not(global_tmr_voter(0)(552));                                                             
                tmr_registers(1)(553)    <= not(global_tmr_voter(1)(552));                                                             
                tmr_registers(2)(553)    <= not(global_tmr_voter(2)(552));                                                             
 
                tmr_registers(0)(554)    <= not(global_tmr_voter(0)(553));                                                             
                tmr_registers(1)(554)    <= not(global_tmr_voter(1)(553));                                                             
                tmr_registers(2)(554)    <= not(global_tmr_voter(2)(553));                                                             
 
                tmr_registers(0)(555)    <= not(global_tmr_voter(0)(554));                                                             
                tmr_registers(1)(555)    <= not(global_tmr_voter(1)(554));                                                             
                tmr_registers(2)(555)    <= not(global_tmr_voter(2)(554));                                                             
 
                tmr_registers(0)(556)    <= not(global_tmr_voter(0)(555));                                                             
                tmr_registers(1)(556)    <= not(global_tmr_voter(1)(555));                                                             
                tmr_registers(2)(556)    <= not(global_tmr_voter(2)(555));                                                             
 
                tmr_registers(0)(557)    <= not(global_tmr_voter(0)(556));                                                             
                tmr_registers(1)(557)    <= not(global_tmr_voter(1)(556));                                                             
                tmr_registers(2)(557)    <= not(global_tmr_voter(2)(556));                                                             
 
                tmr_registers(0)(558)    <= not(global_tmr_voter(0)(557));                                                             
                tmr_registers(1)(558)    <= not(global_tmr_voter(1)(557));                                                             
                tmr_registers(2)(558)    <= not(global_tmr_voter(2)(557));                                                             
 
                tmr_registers(0)(559)    <= not(global_tmr_voter(0)(558));                                                             
                tmr_registers(1)(559)    <= not(global_tmr_voter(1)(558));                                                             
                tmr_registers(2)(559)    <= not(global_tmr_voter(2)(558));                                                             
 
                tmr_registers(0)(560)    <= not(global_tmr_voter(0)(559));                                                             
                tmr_registers(1)(560)    <= not(global_tmr_voter(1)(559));                                                             
                tmr_registers(2)(560)    <= not(global_tmr_voter(2)(559));                                                             
 
                tmr_registers(0)(561)    <= not(global_tmr_voter(0)(560));                                                             
                tmr_registers(1)(561)    <= not(global_tmr_voter(1)(560));                                                             
                tmr_registers(2)(561)    <= not(global_tmr_voter(2)(560));                                                             
 
                tmr_registers(0)(562)    <= not(global_tmr_voter(0)(561));                                                             
                tmr_registers(1)(562)    <= not(global_tmr_voter(1)(561));                                                             
                tmr_registers(2)(562)    <= not(global_tmr_voter(2)(561));                                                             
 
                tmr_registers(0)(563)    <= not(global_tmr_voter(0)(562));                                                             
                tmr_registers(1)(563)    <= not(global_tmr_voter(1)(562));                                                             
                tmr_registers(2)(563)    <= not(global_tmr_voter(2)(562));                                                             
 
                tmr_registers(0)(564)    <= not(global_tmr_voter(0)(563));                                                             
                tmr_registers(1)(564)    <= not(global_tmr_voter(1)(563));                                                             
                tmr_registers(2)(564)    <= not(global_tmr_voter(2)(563));                                                             
 
                tmr_registers(0)(565)    <= not(global_tmr_voter(0)(564));                                                             
                tmr_registers(1)(565)    <= not(global_tmr_voter(1)(564));                                                             
                tmr_registers(2)(565)    <= not(global_tmr_voter(2)(564));                                                             
 
                tmr_registers(0)(566)    <= not(global_tmr_voter(0)(565));                                                             
                tmr_registers(1)(566)    <= not(global_tmr_voter(1)(565));                                                             
                tmr_registers(2)(566)    <= not(global_tmr_voter(2)(565));                                                             
 
                tmr_registers(0)(567)    <= not(global_tmr_voter(0)(566));                                                             
                tmr_registers(1)(567)    <= not(global_tmr_voter(1)(566));                                                             
                tmr_registers(2)(567)    <= not(global_tmr_voter(2)(566));                                                             
 
                tmr_registers(0)(568)    <= not(global_tmr_voter(0)(567));                                                             
                tmr_registers(1)(568)    <= not(global_tmr_voter(1)(567));                                                             
                tmr_registers(2)(568)    <= not(global_tmr_voter(2)(567));                                                             
 
                tmr_registers(0)(569)    <= not(global_tmr_voter(0)(568));                                                             
                tmr_registers(1)(569)    <= not(global_tmr_voter(1)(568));                                                             
                tmr_registers(2)(569)    <= not(global_tmr_voter(2)(568));                                                             
 
                tmr_registers(0)(570)    <= not(global_tmr_voter(0)(569));                                                             
                tmr_registers(1)(570)    <= not(global_tmr_voter(1)(569));                                                             
                tmr_registers(2)(570)    <= not(global_tmr_voter(2)(569));                                                             
 
                tmr_registers(0)(571)    <= not(global_tmr_voter(0)(570));                                                             
                tmr_registers(1)(571)    <= not(global_tmr_voter(1)(570));                                                             
                tmr_registers(2)(571)    <= not(global_tmr_voter(2)(570));                                                             
 
                tmr_registers(0)(572)    <= not(global_tmr_voter(0)(571));                                                             
                tmr_registers(1)(572)    <= not(global_tmr_voter(1)(571));                                                             
                tmr_registers(2)(572)    <= not(global_tmr_voter(2)(571));                                                             
 
                tmr_registers(0)(573)    <= not(global_tmr_voter(0)(572));                                                             
                tmr_registers(1)(573)    <= not(global_tmr_voter(1)(572));                                                             
                tmr_registers(2)(573)    <= not(global_tmr_voter(2)(572));                                                             
 
                tmr_registers(0)(574)    <= not(global_tmr_voter(0)(573));                                                             
                tmr_registers(1)(574)    <= not(global_tmr_voter(1)(573));                                                             
                tmr_registers(2)(574)    <= not(global_tmr_voter(2)(573));                                                             
 
                tmr_registers(0)(575)    <= not(global_tmr_voter(0)(574));                                                             
                tmr_registers(1)(575)    <= not(global_tmr_voter(1)(574));                                                             
                tmr_registers(2)(575)    <= not(global_tmr_voter(2)(574));                                                             
 
                tmr_registers(0)(576)    <= not(global_tmr_voter(0)(575));                                                             
                tmr_registers(1)(576)    <= not(global_tmr_voter(1)(575));                                                             
                tmr_registers(2)(576)    <= not(global_tmr_voter(2)(575));                                                             
 
                tmr_registers(0)(577)    <= not(global_tmr_voter(0)(576));                                                             
                tmr_registers(1)(577)    <= not(global_tmr_voter(1)(576));                                                             
                tmr_registers(2)(577)    <= not(global_tmr_voter(2)(576));                                                             
 
                tmr_registers(0)(578)    <= not(global_tmr_voter(0)(577));                                                             
                tmr_registers(1)(578)    <= not(global_tmr_voter(1)(577));                                                             
                tmr_registers(2)(578)    <= not(global_tmr_voter(2)(577));                                                             
 
                tmr_registers(0)(579)    <= not(global_tmr_voter(0)(578));                                                             
                tmr_registers(1)(579)    <= not(global_tmr_voter(1)(578));                                                             
                tmr_registers(2)(579)    <= not(global_tmr_voter(2)(578));                                                             
 
                tmr_registers(0)(580)    <= not(global_tmr_voter(0)(579));                                                             
                tmr_registers(1)(580)    <= not(global_tmr_voter(1)(579));                                                             
                tmr_registers(2)(580)    <= not(global_tmr_voter(2)(579));                                                             
 
                tmr_registers(0)(581)    <= not(global_tmr_voter(0)(580));                                                             
                tmr_registers(1)(581)    <= not(global_tmr_voter(1)(580));                                                             
                tmr_registers(2)(581)    <= not(global_tmr_voter(2)(580));                                                             
 
                tmr_registers(0)(582)    <= not(global_tmr_voter(0)(581));                                                             
                tmr_registers(1)(582)    <= not(global_tmr_voter(1)(581));                                                             
                tmr_registers(2)(582)    <= not(global_tmr_voter(2)(581));                                                             
 
                tmr_registers(0)(583)    <= not(global_tmr_voter(0)(582));                                                             
                tmr_registers(1)(583)    <= not(global_tmr_voter(1)(582));                                                             
                tmr_registers(2)(583)    <= not(global_tmr_voter(2)(582));                                                             
 
                tmr_registers(0)(584)    <= not(global_tmr_voter(0)(583));                                                             
                tmr_registers(1)(584)    <= not(global_tmr_voter(1)(583));                                                             
                tmr_registers(2)(584)    <= not(global_tmr_voter(2)(583));                                                             
 
                tmr_registers(0)(585)    <= not(global_tmr_voter(0)(584));                                                             
                tmr_registers(1)(585)    <= not(global_tmr_voter(1)(584));                                                             
                tmr_registers(2)(585)    <= not(global_tmr_voter(2)(584));                                                             
 
                tmr_registers(0)(586)    <= not(global_tmr_voter(0)(585));                                                             
                tmr_registers(1)(586)    <= not(global_tmr_voter(1)(585));                                                             
                tmr_registers(2)(586)    <= not(global_tmr_voter(2)(585));                                                             
 
                tmr_registers(0)(587)    <= not(global_tmr_voter(0)(586));                                                             
                tmr_registers(1)(587)    <= not(global_tmr_voter(1)(586));                                                             
                tmr_registers(2)(587)    <= not(global_tmr_voter(2)(586));                                                             
 
                tmr_registers(0)(588)    <= not(global_tmr_voter(0)(587));                                                             
                tmr_registers(1)(588)    <= not(global_tmr_voter(1)(587));                                                             
                tmr_registers(2)(588)    <= not(global_tmr_voter(2)(587));                                                             
 
                tmr_registers(0)(589)    <= not(global_tmr_voter(0)(588));                                                             
                tmr_registers(1)(589)    <= not(global_tmr_voter(1)(588));                                                             
                tmr_registers(2)(589)    <= not(global_tmr_voter(2)(588));                                                             
 
                tmr_registers(0)(590)    <= not(global_tmr_voter(0)(589));                                                             
                tmr_registers(1)(590)    <= not(global_tmr_voter(1)(589));                                                             
                tmr_registers(2)(590)    <= not(global_tmr_voter(2)(589));                                                             
 
                tmr_registers(0)(591)    <= not(global_tmr_voter(0)(590));                                                             
                tmr_registers(1)(591)    <= not(global_tmr_voter(1)(590));                                                             
                tmr_registers(2)(591)    <= not(global_tmr_voter(2)(590));                                                             
 
                tmr_registers(0)(592)    <= not(global_tmr_voter(0)(591));                                                             
                tmr_registers(1)(592)    <= not(global_tmr_voter(1)(591));                                                             
                tmr_registers(2)(592)    <= not(global_tmr_voter(2)(591));                                                             
 
                tmr_registers(0)(593)    <= not(global_tmr_voter(0)(592));                                                             
                tmr_registers(1)(593)    <= not(global_tmr_voter(1)(592));                                                             
                tmr_registers(2)(593)    <= not(global_tmr_voter(2)(592));                                                             
 
                tmr_registers(0)(594)    <= not(global_tmr_voter(0)(593));                                                             
                tmr_registers(1)(594)    <= not(global_tmr_voter(1)(593));                                                             
                tmr_registers(2)(594)    <= not(global_tmr_voter(2)(593));                                                             
 
                tmr_registers(0)(595)    <= not(global_tmr_voter(0)(594));                                                             
                tmr_registers(1)(595)    <= not(global_tmr_voter(1)(594));                                                             
                tmr_registers(2)(595)    <= not(global_tmr_voter(2)(594));                                                             
 
                tmr_registers(0)(596)    <= not(global_tmr_voter(0)(595));                                                             
                tmr_registers(1)(596)    <= not(global_tmr_voter(1)(595));                                                             
                tmr_registers(2)(596)    <= not(global_tmr_voter(2)(595));                                                             
 
                tmr_registers(0)(597)    <= not(global_tmr_voter(0)(596));                                                             
                tmr_registers(1)(597)    <= not(global_tmr_voter(1)(596));                                                             
                tmr_registers(2)(597)    <= not(global_tmr_voter(2)(596));                                                             
 
                tmr_registers(0)(598)    <= not(global_tmr_voter(0)(597));                                                             
                tmr_registers(1)(598)    <= not(global_tmr_voter(1)(597));                                                             
                tmr_registers(2)(598)    <= not(global_tmr_voter(2)(597));                                                             
 
                tmr_registers(0)(599)    <= not(global_tmr_voter(0)(598));                                                             
                tmr_registers(1)(599)    <= not(global_tmr_voter(1)(598));                                                             
                tmr_registers(2)(599)    <= not(global_tmr_voter(2)(598));                                                             
 
                tmr_registers(0)(600)    <= not(global_tmr_voter(0)(599));                                                             
                tmr_registers(1)(600)    <= not(global_tmr_voter(1)(599));                                                             
                tmr_registers(2)(600)    <= not(global_tmr_voter(2)(599));                                                             
 
                tmr_registers(0)(601)    <= not(global_tmr_voter(0)(600));                                                             
                tmr_registers(1)(601)    <= not(global_tmr_voter(1)(600));                                                             
                tmr_registers(2)(601)    <= not(global_tmr_voter(2)(600));                                                             
 
                tmr_registers(0)(602)    <= not(global_tmr_voter(0)(601));                                                             
                tmr_registers(1)(602)    <= not(global_tmr_voter(1)(601));                                                             
                tmr_registers(2)(602)    <= not(global_tmr_voter(2)(601));                                                             
 
                tmr_registers(0)(603)    <= not(global_tmr_voter(0)(602));                                                             
                tmr_registers(1)(603)    <= not(global_tmr_voter(1)(602));                                                             
                tmr_registers(2)(603)    <= not(global_tmr_voter(2)(602));                                                             
 
                tmr_registers(0)(604)    <= not(global_tmr_voter(0)(603));                                                             
                tmr_registers(1)(604)    <= not(global_tmr_voter(1)(603));                                                             
                tmr_registers(2)(604)    <= not(global_tmr_voter(2)(603));                                                             
 
                tmr_registers(0)(605)    <= not(global_tmr_voter(0)(604));                                                             
                tmr_registers(1)(605)    <= not(global_tmr_voter(1)(604));                                                             
                tmr_registers(2)(605)    <= not(global_tmr_voter(2)(604));                                                             
 
                tmr_registers(0)(606)    <= not(global_tmr_voter(0)(605));                                                             
                tmr_registers(1)(606)    <= not(global_tmr_voter(1)(605));                                                             
                tmr_registers(2)(606)    <= not(global_tmr_voter(2)(605));                                                             
 
                tmr_registers(0)(607)    <= not(global_tmr_voter(0)(606));                                                             
                tmr_registers(1)(607)    <= not(global_tmr_voter(1)(606));                                                             
                tmr_registers(2)(607)    <= not(global_tmr_voter(2)(606));                                                             
 
                tmr_registers(0)(608)    <= not(global_tmr_voter(0)(607));                                                             
                tmr_registers(1)(608)    <= not(global_tmr_voter(1)(607));                                                             
                tmr_registers(2)(608)    <= not(global_tmr_voter(2)(607));                                                             
 
                tmr_registers(0)(609)    <= not(global_tmr_voter(0)(608));                                                             
                tmr_registers(1)(609)    <= not(global_tmr_voter(1)(608));                                                             
                tmr_registers(2)(609)    <= not(global_tmr_voter(2)(608));                                                             
 
                tmr_registers(0)(610)    <= not(global_tmr_voter(0)(609));                                                             
                tmr_registers(1)(610)    <= not(global_tmr_voter(1)(609));                                                             
                tmr_registers(2)(610)    <= not(global_tmr_voter(2)(609));                                                             
 
                tmr_registers(0)(611)    <= not(global_tmr_voter(0)(610));                                                             
                tmr_registers(1)(611)    <= not(global_tmr_voter(1)(610));                                                             
                tmr_registers(2)(611)    <= not(global_tmr_voter(2)(610));                                                             
 
                tmr_registers(0)(612)    <= not(global_tmr_voter(0)(611));                                                             
                tmr_registers(1)(612)    <= not(global_tmr_voter(1)(611));                                                             
                tmr_registers(2)(612)    <= not(global_tmr_voter(2)(611));                                                             
 
                tmr_registers(0)(613)    <= not(global_tmr_voter(0)(612));                                                             
                tmr_registers(1)(613)    <= not(global_tmr_voter(1)(612));                                                             
                tmr_registers(2)(613)    <= not(global_tmr_voter(2)(612));                                                             
 
                tmr_registers(0)(614)    <= not(global_tmr_voter(0)(613));                                                             
                tmr_registers(1)(614)    <= not(global_tmr_voter(1)(613));                                                             
                tmr_registers(2)(614)    <= not(global_tmr_voter(2)(613));                                                             
 
                tmr_registers(0)(615)    <= not(global_tmr_voter(0)(614));                                                             
                tmr_registers(1)(615)    <= not(global_tmr_voter(1)(614));                                                             
                tmr_registers(2)(615)    <= not(global_tmr_voter(2)(614));                                                             
 
                tmr_registers(0)(616)    <= not(global_tmr_voter(0)(615));                                                             
                tmr_registers(1)(616)    <= not(global_tmr_voter(1)(615));                                                             
                tmr_registers(2)(616)    <= not(global_tmr_voter(2)(615));                                                             
 
                tmr_registers(0)(617)    <= not(global_tmr_voter(0)(616));                                                             
                tmr_registers(1)(617)    <= not(global_tmr_voter(1)(616));                                                             
                tmr_registers(2)(617)    <= not(global_tmr_voter(2)(616));                                                             
 
                tmr_registers(0)(618)    <= not(global_tmr_voter(0)(617));                                                             
                tmr_registers(1)(618)    <= not(global_tmr_voter(1)(617));                                                             
                tmr_registers(2)(618)    <= not(global_tmr_voter(2)(617));                                                             
 
                tmr_registers(0)(619)    <= not(global_tmr_voter(0)(618));                                                             
                tmr_registers(1)(619)    <= not(global_tmr_voter(1)(618));                                                             
                tmr_registers(2)(619)    <= not(global_tmr_voter(2)(618));                                                             
 
                tmr_registers(0)(620)    <= not(global_tmr_voter(0)(619));                                                             
                tmr_registers(1)(620)    <= not(global_tmr_voter(1)(619));                                                             
                tmr_registers(2)(620)    <= not(global_tmr_voter(2)(619));                                                             
 
                tmr_registers(0)(621)    <= not(global_tmr_voter(0)(620));                                                             
                tmr_registers(1)(621)    <= not(global_tmr_voter(1)(620));                                                             
                tmr_registers(2)(621)    <= not(global_tmr_voter(2)(620));                                                             
 
                tmr_registers(0)(622)    <= not(global_tmr_voter(0)(621));                                                             
                tmr_registers(1)(622)    <= not(global_tmr_voter(1)(621));                                                             
                tmr_registers(2)(622)    <= not(global_tmr_voter(2)(621));                                                             
 
                tmr_registers(0)(623)    <= not(global_tmr_voter(0)(622));                                                             
                tmr_registers(1)(623)    <= not(global_tmr_voter(1)(622));                                                             
                tmr_registers(2)(623)    <= not(global_tmr_voter(2)(622));                                                             
 
                tmr_registers(0)(624)    <= not(global_tmr_voter(0)(623));                                                             
                tmr_registers(1)(624)    <= not(global_tmr_voter(1)(623));                                                             
                tmr_registers(2)(624)    <= not(global_tmr_voter(2)(623));                                                             
 
                tmr_registers(0)(625)    <= not(global_tmr_voter(0)(624));                                                             
                tmr_registers(1)(625)    <= not(global_tmr_voter(1)(624));                                                             
                tmr_registers(2)(625)    <= not(global_tmr_voter(2)(624));                                                             
 
                tmr_registers(0)(626)    <= not(global_tmr_voter(0)(625));                                                             
                tmr_registers(1)(626)    <= not(global_tmr_voter(1)(625));                                                             
                tmr_registers(2)(626)    <= not(global_tmr_voter(2)(625));                                                             
 
                tmr_registers(0)(627)    <= not(global_tmr_voter(0)(626));                                                             
                tmr_registers(1)(627)    <= not(global_tmr_voter(1)(626));                                                             
                tmr_registers(2)(627)    <= not(global_tmr_voter(2)(626));                                                             
 
                tmr_registers(0)(628)    <= not(global_tmr_voter(0)(627));                                                             
                tmr_registers(1)(628)    <= not(global_tmr_voter(1)(627));                                                             
                tmr_registers(2)(628)    <= not(global_tmr_voter(2)(627));                                                             
 
                tmr_registers(0)(629)    <= not(global_tmr_voter(0)(628));                                                             
                tmr_registers(1)(629)    <= not(global_tmr_voter(1)(628));                                                             
                tmr_registers(2)(629)    <= not(global_tmr_voter(2)(628));                                                             
 
                tmr_registers(0)(630)    <= not(global_tmr_voter(0)(629));                                                             
                tmr_registers(1)(630)    <= not(global_tmr_voter(1)(629));                                                             
                tmr_registers(2)(630)    <= not(global_tmr_voter(2)(629));                                                             
 
                tmr_registers(0)(631)    <= not(global_tmr_voter(0)(630));                                                             
                tmr_registers(1)(631)    <= not(global_tmr_voter(1)(630));                                                             
                tmr_registers(2)(631)    <= not(global_tmr_voter(2)(630));                                                             
 
                tmr_registers(0)(632)    <= not(global_tmr_voter(0)(631));                                                             
                tmr_registers(1)(632)    <= not(global_tmr_voter(1)(631));                                                             
                tmr_registers(2)(632)    <= not(global_tmr_voter(2)(631));                                                             
 
                tmr_registers(0)(633)    <= not(global_tmr_voter(0)(632));                                                             
                tmr_registers(1)(633)    <= not(global_tmr_voter(1)(632));                                                             
                tmr_registers(2)(633)    <= not(global_tmr_voter(2)(632));                                                             
 
                tmr_registers(0)(634)    <= not(global_tmr_voter(0)(633));                                                             
                tmr_registers(1)(634)    <= not(global_tmr_voter(1)(633));                                                             
                tmr_registers(2)(634)    <= not(global_tmr_voter(2)(633));                                                             
 
                tmr_registers(0)(635)    <= not(global_tmr_voter(0)(634));                                                             
                tmr_registers(1)(635)    <= not(global_tmr_voter(1)(634));                                                             
                tmr_registers(2)(635)    <= not(global_tmr_voter(2)(634));                                                             
 
                tmr_registers(0)(636)    <= not(global_tmr_voter(0)(635));                                                             
                tmr_registers(1)(636)    <= not(global_tmr_voter(1)(635));                                                             
                tmr_registers(2)(636)    <= not(global_tmr_voter(2)(635));                                                             
 
                tmr_registers(0)(637)    <= not(global_tmr_voter(0)(636));                                                             
                tmr_registers(1)(637)    <= not(global_tmr_voter(1)(636));                                                             
                tmr_registers(2)(637)    <= not(global_tmr_voter(2)(636));                                                             
 
                tmr_registers(0)(638)    <= not(global_tmr_voter(0)(637));                                                             
                tmr_registers(1)(638)    <= not(global_tmr_voter(1)(637));                                                             
                tmr_registers(2)(638)    <= not(global_tmr_voter(2)(637));                                                             
 
                tmr_registers(0)(639)    <= not(global_tmr_voter(0)(638));                                                             
                tmr_registers(1)(639)    <= not(global_tmr_voter(1)(638));                                                             
                tmr_registers(2)(639)    <= not(global_tmr_voter(2)(638));                                                             
 
                tmr_registers(0)(640)    <= not(global_tmr_voter(0)(639));                                                             
                tmr_registers(1)(640)    <= not(global_tmr_voter(1)(639));                                                             
                tmr_registers(2)(640)    <= not(global_tmr_voter(2)(639));                                                             
 
                tmr_registers(0)(641)    <= not(global_tmr_voter(0)(640));                                                             
                tmr_registers(1)(641)    <= not(global_tmr_voter(1)(640));                                                             
                tmr_registers(2)(641)    <= not(global_tmr_voter(2)(640));                                                             
 
                tmr_registers(0)(642)    <= not(global_tmr_voter(0)(641));                                                             
                tmr_registers(1)(642)    <= not(global_tmr_voter(1)(641));                                                             
                tmr_registers(2)(642)    <= not(global_tmr_voter(2)(641));                                                             
 
                tmr_registers(0)(643)    <= not(global_tmr_voter(0)(642));                                                             
                tmr_registers(1)(643)    <= not(global_tmr_voter(1)(642));                                                             
                tmr_registers(2)(643)    <= not(global_tmr_voter(2)(642));                                                             
 
                tmr_registers(0)(644)    <= not(global_tmr_voter(0)(643));                                                             
                tmr_registers(1)(644)    <= not(global_tmr_voter(1)(643));                                                             
                tmr_registers(2)(644)    <= not(global_tmr_voter(2)(643));                                                             
 
                tmr_registers(0)(645)    <= not(global_tmr_voter(0)(644));                                                             
                tmr_registers(1)(645)    <= not(global_tmr_voter(1)(644));                                                             
                tmr_registers(2)(645)    <= not(global_tmr_voter(2)(644));                                                             
 
                tmr_registers(0)(646)    <= not(global_tmr_voter(0)(645));                                                             
                tmr_registers(1)(646)    <= not(global_tmr_voter(1)(645));                                                             
                tmr_registers(2)(646)    <= not(global_tmr_voter(2)(645));                                                             
 
                tmr_registers(0)(647)    <= not(global_tmr_voter(0)(646));                                                             
                tmr_registers(1)(647)    <= not(global_tmr_voter(1)(646));                                                             
                tmr_registers(2)(647)    <= not(global_tmr_voter(2)(646));                                                             
 
                tmr_registers(0)(648)    <= not(global_tmr_voter(0)(647));                                                             
                tmr_registers(1)(648)    <= not(global_tmr_voter(1)(647));                                                             
                tmr_registers(2)(648)    <= not(global_tmr_voter(2)(647));                                                             
 
                tmr_registers(0)(649)    <= not(global_tmr_voter(0)(648));                                                             
                tmr_registers(1)(649)    <= not(global_tmr_voter(1)(648));                                                             
                tmr_registers(2)(649)    <= not(global_tmr_voter(2)(648));                                                             
 
                tmr_registers(0)(650)    <= not(global_tmr_voter(0)(649));                                                             
                tmr_registers(1)(650)    <= not(global_tmr_voter(1)(649));                                                             
                tmr_registers(2)(650)    <= not(global_tmr_voter(2)(649));                                                             
 
                tmr_registers(0)(651)    <= not(global_tmr_voter(0)(650));                                                             
                tmr_registers(1)(651)    <= not(global_tmr_voter(1)(650));                                                             
                tmr_registers(2)(651)    <= not(global_tmr_voter(2)(650));                                                             
 
                tmr_registers(0)(652)    <= not(global_tmr_voter(0)(651));                                                             
                tmr_registers(1)(652)    <= not(global_tmr_voter(1)(651));                                                             
                tmr_registers(2)(652)    <= not(global_tmr_voter(2)(651));                                                             
 
                tmr_registers(0)(653)    <= not(global_tmr_voter(0)(652));                                                             
                tmr_registers(1)(653)    <= not(global_tmr_voter(1)(652));                                                             
                tmr_registers(2)(653)    <= not(global_tmr_voter(2)(652));                                                             
 
                tmr_registers(0)(654)    <= not(global_tmr_voter(0)(653));                                                             
                tmr_registers(1)(654)    <= not(global_tmr_voter(1)(653));                                                             
                tmr_registers(2)(654)    <= not(global_tmr_voter(2)(653));                                                             
 
                tmr_registers(0)(655)    <= not(global_tmr_voter(0)(654));                                                             
                tmr_registers(1)(655)    <= not(global_tmr_voter(1)(654));                                                             
                tmr_registers(2)(655)    <= not(global_tmr_voter(2)(654));                                                             
 
                tmr_registers(0)(656)    <= not(global_tmr_voter(0)(655));                                                             
                tmr_registers(1)(656)    <= not(global_tmr_voter(1)(655));                                                             
                tmr_registers(2)(656)    <= not(global_tmr_voter(2)(655));                                                             
 
                tmr_registers(0)(657)    <= not(global_tmr_voter(0)(656));                                                             
                tmr_registers(1)(657)    <= not(global_tmr_voter(1)(656));                                                             
                tmr_registers(2)(657)    <= not(global_tmr_voter(2)(656));                                                             
 
                tmr_registers(0)(658)    <= not(global_tmr_voter(0)(657));                                                             
                tmr_registers(1)(658)    <= not(global_tmr_voter(1)(657));                                                             
                tmr_registers(2)(658)    <= not(global_tmr_voter(2)(657));                                                             
 
                tmr_registers(0)(659)    <= not(global_tmr_voter(0)(658));                                                             
                tmr_registers(1)(659)    <= not(global_tmr_voter(1)(658));                                                             
                tmr_registers(2)(659)    <= not(global_tmr_voter(2)(658));                                                             
 
                tmr_registers(0)(660)    <= not(global_tmr_voter(0)(659));                                                             
                tmr_registers(1)(660)    <= not(global_tmr_voter(1)(659));                                                             
                tmr_registers(2)(660)    <= not(global_tmr_voter(2)(659));                                                             
 
                tmr_registers(0)(661)    <= not(global_tmr_voter(0)(660));                                                             
                tmr_registers(1)(661)    <= not(global_tmr_voter(1)(660));                                                             
                tmr_registers(2)(661)    <= not(global_tmr_voter(2)(660));                                                             
 
                tmr_registers(0)(662)    <= not(global_tmr_voter(0)(661));                                                             
                tmr_registers(1)(662)    <= not(global_tmr_voter(1)(661));                                                             
                tmr_registers(2)(662)    <= not(global_tmr_voter(2)(661));                                                             
 
                tmr_registers(0)(663)    <= not(global_tmr_voter(0)(662));                                                             
                tmr_registers(1)(663)    <= not(global_tmr_voter(1)(662));                                                             
                tmr_registers(2)(663)    <= not(global_tmr_voter(2)(662));                                                             
 
                tmr_registers(0)(664)    <= not(global_tmr_voter(0)(663));                                                             
                tmr_registers(1)(664)    <= not(global_tmr_voter(1)(663));                                                             
                tmr_registers(2)(664)    <= not(global_tmr_voter(2)(663));                                                             
 
                tmr_registers(0)(665)    <= not(global_tmr_voter(0)(664));                                                             
                tmr_registers(1)(665)    <= not(global_tmr_voter(1)(664));                                                             
                tmr_registers(2)(665)    <= not(global_tmr_voter(2)(664));                                                             
 
                tmr_registers(0)(666)    <= not(global_tmr_voter(0)(665));                                                             
                tmr_registers(1)(666)    <= not(global_tmr_voter(1)(665));                                                             
                tmr_registers(2)(666)    <= not(global_tmr_voter(2)(665));                                                             
 
                tmr_registers(0)(667)    <= not(global_tmr_voter(0)(666));                                                             
                tmr_registers(1)(667)    <= not(global_tmr_voter(1)(666));                                                             
                tmr_registers(2)(667)    <= not(global_tmr_voter(2)(666));                                                             
 
                tmr_registers(0)(668)    <= not(global_tmr_voter(0)(667));                                                             
                tmr_registers(1)(668)    <= not(global_tmr_voter(1)(667));                                                             
                tmr_registers(2)(668)    <= not(global_tmr_voter(2)(667));                                                             
 
                tmr_registers(0)(669)    <= not(global_tmr_voter(0)(668));                                                             
                tmr_registers(1)(669)    <= not(global_tmr_voter(1)(668));                                                             
                tmr_registers(2)(669)    <= not(global_tmr_voter(2)(668));                                                             
 
                tmr_registers(0)(670)    <= not(global_tmr_voter(0)(669));                                                             
                tmr_registers(1)(670)    <= not(global_tmr_voter(1)(669));                                                             
                tmr_registers(2)(670)    <= not(global_tmr_voter(2)(669));                                                             
 
                tmr_registers(0)(671)    <= not(global_tmr_voter(0)(670));                                                             
                tmr_registers(1)(671)    <= not(global_tmr_voter(1)(670));                                                             
                tmr_registers(2)(671)    <= not(global_tmr_voter(2)(670));                                                             
 
                tmr_registers(0)(672)    <= not(global_tmr_voter(0)(671));                                                             
                tmr_registers(1)(672)    <= not(global_tmr_voter(1)(671));                                                             
                tmr_registers(2)(672)    <= not(global_tmr_voter(2)(671));                                                             
 
                tmr_registers(0)(673)    <= not(global_tmr_voter(0)(672));                                                             
                tmr_registers(1)(673)    <= not(global_tmr_voter(1)(672));                                                             
                tmr_registers(2)(673)    <= not(global_tmr_voter(2)(672));                                                             
 
                tmr_registers(0)(674)    <= not(global_tmr_voter(0)(673));                                                             
                tmr_registers(1)(674)    <= not(global_tmr_voter(1)(673));                                                             
                tmr_registers(2)(674)    <= not(global_tmr_voter(2)(673));                                                             
 
                tmr_registers(0)(675)    <= not(global_tmr_voter(0)(674));                                                             
                tmr_registers(1)(675)    <= not(global_tmr_voter(1)(674));                                                             
                tmr_registers(2)(675)    <= not(global_tmr_voter(2)(674));                                                             
 
                tmr_registers(0)(676)    <= not(global_tmr_voter(0)(675));                                                             
                tmr_registers(1)(676)    <= not(global_tmr_voter(1)(675));                                                             
                tmr_registers(2)(676)    <= not(global_tmr_voter(2)(675));                                                             
 
                tmr_registers(0)(677)    <= not(global_tmr_voter(0)(676));                                                             
                tmr_registers(1)(677)    <= not(global_tmr_voter(1)(676));                                                             
                tmr_registers(2)(677)    <= not(global_tmr_voter(2)(676));                                                             
 
                tmr_registers(0)(678)    <= not(global_tmr_voter(0)(677));                                                             
                tmr_registers(1)(678)    <= not(global_tmr_voter(1)(677));                                                             
                tmr_registers(2)(678)    <= not(global_tmr_voter(2)(677));                                                             
 
                tmr_registers(0)(679)    <= not(global_tmr_voter(0)(678));                                                             
                tmr_registers(1)(679)    <= not(global_tmr_voter(1)(678));                                                             
                tmr_registers(2)(679)    <= not(global_tmr_voter(2)(678));                                                             
 
                tmr_registers(0)(680)    <= not(global_tmr_voter(0)(679));                                                             
                tmr_registers(1)(680)    <= not(global_tmr_voter(1)(679));                                                             
                tmr_registers(2)(680)    <= not(global_tmr_voter(2)(679));                                                             
 
                tmr_registers(0)(681)    <= not(global_tmr_voter(0)(680));                                                             
                tmr_registers(1)(681)    <= not(global_tmr_voter(1)(680));                                                             
                tmr_registers(2)(681)    <= not(global_tmr_voter(2)(680));                                                             
 
                tmr_registers(0)(682)    <= not(global_tmr_voter(0)(681));                                                             
                tmr_registers(1)(682)    <= not(global_tmr_voter(1)(681));                                                             
                tmr_registers(2)(682)    <= not(global_tmr_voter(2)(681));                                                             
 
                tmr_registers(0)(683)    <= not(global_tmr_voter(0)(682));                                                             
                tmr_registers(1)(683)    <= not(global_tmr_voter(1)(682));                                                             
                tmr_registers(2)(683)    <= not(global_tmr_voter(2)(682));                                                             
 
                tmr_registers(0)(684)    <= not(global_tmr_voter(0)(683));                                                             
                tmr_registers(1)(684)    <= not(global_tmr_voter(1)(683));                                                             
                tmr_registers(2)(684)    <= not(global_tmr_voter(2)(683));                                                             
 
                tmr_registers(0)(685)    <= not(global_tmr_voter(0)(684));                                                             
                tmr_registers(1)(685)    <= not(global_tmr_voter(1)(684));                                                             
                tmr_registers(2)(685)    <= not(global_tmr_voter(2)(684));                                                             
 
                tmr_registers(0)(686)    <= not(global_tmr_voter(0)(685));                                                             
                tmr_registers(1)(686)    <= not(global_tmr_voter(1)(685));                                                             
                tmr_registers(2)(686)    <= not(global_tmr_voter(2)(685));                                                             
 
                tmr_registers(0)(687)    <= not(global_tmr_voter(0)(686));                                                             
                tmr_registers(1)(687)    <= not(global_tmr_voter(1)(686));                                                             
                tmr_registers(2)(687)    <= not(global_tmr_voter(2)(686));                                                             
 
                tmr_registers(0)(688)    <= not(global_tmr_voter(0)(687));                                                             
                tmr_registers(1)(688)    <= not(global_tmr_voter(1)(687));                                                             
                tmr_registers(2)(688)    <= not(global_tmr_voter(2)(687));                                                             
 
                tmr_registers(0)(689)    <= not(global_tmr_voter(0)(688));                                                             
                tmr_registers(1)(689)    <= not(global_tmr_voter(1)(688));                                                             
                tmr_registers(2)(689)    <= not(global_tmr_voter(2)(688));                                                             
 
                tmr_registers(0)(690)    <= not(global_tmr_voter(0)(689));                                                             
                tmr_registers(1)(690)    <= not(global_tmr_voter(1)(689));                                                             
                tmr_registers(2)(690)    <= not(global_tmr_voter(2)(689));                                                             
 
                tmr_registers(0)(691)    <= not(global_tmr_voter(0)(690));                                                             
                tmr_registers(1)(691)    <= not(global_tmr_voter(1)(690));                                                             
                tmr_registers(2)(691)    <= not(global_tmr_voter(2)(690));                                                             
 
                tmr_registers(0)(692)    <= not(global_tmr_voter(0)(691));                                                             
                tmr_registers(1)(692)    <= not(global_tmr_voter(1)(691));                                                             
                tmr_registers(2)(692)    <= not(global_tmr_voter(2)(691));                                                             
 
                tmr_registers(0)(693)    <= not(global_tmr_voter(0)(692));                                                             
                tmr_registers(1)(693)    <= not(global_tmr_voter(1)(692));                                                             
                tmr_registers(2)(693)    <= not(global_tmr_voter(2)(692));                                                             
 
                tmr_registers(0)(694)    <= not(global_tmr_voter(0)(693));                                                             
                tmr_registers(1)(694)    <= not(global_tmr_voter(1)(693));                                                             
                tmr_registers(2)(694)    <= not(global_tmr_voter(2)(693));                                                             
 
                tmr_registers(0)(695)    <= not(global_tmr_voter(0)(694));                                                             
                tmr_registers(1)(695)    <= not(global_tmr_voter(1)(694));                                                             
                tmr_registers(2)(695)    <= not(global_tmr_voter(2)(694));                                                             
 
                tmr_registers(0)(696)    <= not(global_tmr_voter(0)(695));                                                             
                tmr_registers(1)(696)    <= not(global_tmr_voter(1)(695));                                                             
                tmr_registers(2)(696)    <= not(global_tmr_voter(2)(695));                                                             
 
                tmr_registers(0)(697)    <= not(global_tmr_voter(0)(696));                                                             
                tmr_registers(1)(697)    <= not(global_tmr_voter(1)(696));                                                             
                tmr_registers(2)(697)    <= not(global_tmr_voter(2)(696));                                                             
 
                tmr_registers(0)(698)    <= not(global_tmr_voter(0)(697));                                                             
                tmr_registers(1)(698)    <= not(global_tmr_voter(1)(697));                                                             
                tmr_registers(2)(698)    <= not(global_tmr_voter(2)(697));                                                             
 
                tmr_registers(0)(699)    <= not(global_tmr_voter(0)(698));                                                             
                tmr_registers(1)(699)    <= not(global_tmr_voter(1)(698));                                                             
                tmr_registers(2)(699)    <= not(global_tmr_voter(2)(698));                                                             
 
                tmr_registers(0)(700)    <= not(global_tmr_voter(0)(699));                                                             
                tmr_registers(1)(700)    <= not(global_tmr_voter(1)(699));                                                             
                tmr_registers(2)(700)    <= not(global_tmr_voter(2)(699));                                                             
 
                tmr_registers(0)(701)    <= not(global_tmr_voter(0)(700));                                                             
                tmr_registers(1)(701)    <= not(global_tmr_voter(1)(700));                                                             
                tmr_registers(2)(701)    <= not(global_tmr_voter(2)(700));                                                             
 
                tmr_registers(0)(702)    <= not(global_tmr_voter(0)(701));                                                             
                tmr_registers(1)(702)    <= not(global_tmr_voter(1)(701));                                                             
                tmr_registers(2)(702)    <= not(global_tmr_voter(2)(701));                                                             
 
                tmr_registers(0)(703)    <= not(global_tmr_voter(0)(702));                                                             
                tmr_registers(1)(703)    <= not(global_tmr_voter(1)(702));                                                             
                tmr_registers(2)(703)    <= not(global_tmr_voter(2)(702));                                                             
 
                tmr_registers(0)(704)    <= not(global_tmr_voter(0)(703));                                                             
                tmr_registers(1)(704)    <= not(global_tmr_voter(1)(703));                                                             
                tmr_registers(2)(704)    <= not(global_tmr_voter(2)(703));                                                             
 
                tmr_registers(0)(705)    <= not(global_tmr_voter(0)(704));                                                             
                tmr_registers(1)(705)    <= not(global_tmr_voter(1)(704));                                                             
                tmr_registers(2)(705)    <= not(global_tmr_voter(2)(704));                                                             
 
                tmr_registers(0)(706)    <= not(global_tmr_voter(0)(705));                                                             
                tmr_registers(1)(706)    <= not(global_tmr_voter(1)(705));                                                             
                tmr_registers(2)(706)    <= not(global_tmr_voter(2)(705));                                                             
 
                tmr_registers(0)(707)    <= not(global_tmr_voter(0)(706));                                                             
                tmr_registers(1)(707)    <= not(global_tmr_voter(1)(706));                                                             
                tmr_registers(2)(707)    <= not(global_tmr_voter(2)(706));                                                             
 
                tmr_registers(0)(708)    <= not(global_tmr_voter(0)(707));                                                             
                tmr_registers(1)(708)    <= not(global_tmr_voter(1)(707));                                                             
                tmr_registers(2)(708)    <= not(global_tmr_voter(2)(707));                                                             
 
                tmr_registers(0)(709)    <= not(global_tmr_voter(0)(708));                                                             
                tmr_registers(1)(709)    <= not(global_tmr_voter(1)(708));                                                             
                tmr_registers(2)(709)    <= not(global_tmr_voter(2)(708));                                                             
 
                tmr_registers(0)(710)    <= not(global_tmr_voter(0)(709));                                                             
                tmr_registers(1)(710)    <= not(global_tmr_voter(1)(709));                                                             
                tmr_registers(2)(710)    <= not(global_tmr_voter(2)(709));                                                             
 
                tmr_registers(0)(711)    <= not(global_tmr_voter(0)(710));                                                             
                tmr_registers(1)(711)    <= not(global_tmr_voter(1)(710));                                                             
                tmr_registers(2)(711)    <= not(global_tmr_voter(2)(710));                                                             
 
                tmr_registers(0)(712)    <= not(global_tmr_voter(0)(711));                                                             
                tmr_registers(1)(712)    <= not(global_tmr_voter(1)(711));                                                             
                tmr_registers(2)(712)    <= not(global_tmr_voter(2)(711));                                                             
 
                tmr_registers(0)(713)    <= not(global_tmr_voter(0)(712));                                                             
                tmr_registers(1)(713)    <= not(global_tmr_voter(1)(712));                                                             
                tmr_registers(2)(713)    <= not(global_tmr_voter(2)(712));                                                             
 
                tmr_registers(0)(714)    <= not(global_tmr_voter(0)(713));                                                             
                tmr_registers(1)(714)    <= not(global_tmr_voter(1)(713));                                                             
                tmr_registers(2)(714)    <= not(global_tmr_voter(2)(713));                                                             
 
                tmr_registers(0)(715)    <= not(global_tmr_voter(0)(714));                                                             
                tmr_registers(1)(715)    <= not(global_tmr_voter(1)(714));                                                             
                tmr_registers(2)(715)    <= not(global_tmr_voter(2)(714));                                                             
 
                tmr_registers(0)(716)    <= not(global_tmr_voter(0)(715));                                                             
                tmr_registers(1)(716)    <= not(global_tmr_voter(1)(715));                                                             
                tmr_registers(2)(716)    <= not(global_tmr_voter(2)(715));                                                             
 
                tmr_registers(0)(717)    <= not(global_tmr_voter(0)(716));                                                             
                tmr_registers(1)(717)    <= not(global_tmr_voter(1)(716));                                                             
                tmr_registers(2)(717)    <= not(global_tmr_voter(2)(716));                                                             
 
                tmr_registers(0)(718)    <= not(global_tmr_voter(0)(717));                                                             
                tmr_registers(1)(718)    <= not(global_tmr_voter(1)(717));                                                             
                tmr_registers(2)(718)    <= not(global_tmr_voter(2)(717));                                                             
 
                tmr_registers(0)(719)    <= not(global_tmr_voter(0)(718));                                                             
                tmr_registers(1)(719)    <= not(global_tmr_voter(1)(718));                                                             
                tmr_registers(2)(719)    <= not(global_tmr_voter(2)(718));                                                             
 
                tmr_registers(0)(720)    <= not(global_tmr_voter(0)(719));                                                             
                tmr_registers(1)(720)    <= not(global_tmr_voter(1)(719));                                                             
                tmr_registers(2)(720)    <= not(global_tmr_voter(2)(719));                                                             
 
                tmr_registers(0)(721)    <= not(global_tmr_voter(0)(720));                                                             
                tmr_registers(1)(721)    <= not(global_tmr_voter(1)(720));                                                             
                tmr_registers(2)(721)    <= not(global_tmr_voter(2)(720));                                                             
 
                tmr_registers(0)(722)    <= not(global_tmr_voter(0)(721));                                                             
                tmr_registers(1)(722)    <= not(global_tmr_voter(1)(721));                                                             
                tmr_registers(2)(722)    <= not(global_tmr_voter(2)(721));                                                             
 
                tmr_registers(0)(723)    <= not(global_tmr_voter(0)(722));                                                             
                tmr_registers(1)(723)    <= not(global_tmr_voter(1)(722));                                                             
                tmr_registers(2)(723)    <= not(global_tmr_voter(2)(722));                                                             
 
                tmr_registers(0)(724)    <= not(global_tmr_voter(0)(723));                                                             
                tmr_registers(1)(724)    <= not(global_tmr_voter(1)(723));                                                             
                tmr_registers(2)(724)    <= not(global_tmr_voter(2)(723));                                                             
 
                tmr_registers(0)(725)    <= not(global_tmr_voter(0)(724));                                                             
                tmr_registers(1)(725)    <= not(global_tmr_voter(1)(724));                                                             
                tmr_registers(2)(725)    <= not(global_tmr_voter(2)(724));                                                             
 
                tmr_registers(0)(726)    <= not(global_tmr_voter(0)(725));                                                             
                tmr_registers(1)(726)    <= not(global_tmr_voter(1)(725));                                                             
                tmr_registers(2)(726)    <= not(global_tmr_voter(2)(725));                                                             
 
                tmr_registers(0)(727)    <= not(global_tmr_voter(0)(726));                                                             
                tmr_registers(1)(727)    <= not(global_tmr_voter(1)(726));                                                             
                tmr_registers(2)(727)    <= not(global_tmr_voter(2)(726));                                                             
 
                tmr_registers(0)(728)    <= not(global_tmr_voter(0)(727));                                                             
                tmr_registers(1)(728)    <= not(global_tmr_voter(1)(727));                                                             
                tmr_registers(2)(728)    <= not(global_tmr_voter(2)(727));                                                             
 
                tmr_registers(0)(729)    <= not(global_tmr_voter(0)(728));                                                             
                tmr_registers(1)(729)    <= not(global_tmr_voter(1)(728));                                                             
                tmr_registers(2)(729)    <= not(global_tmr_voter(2)(728));                                                             
 
                tmr_registers(0)(730)    <= not(global_tmr_voter(0)(729));                                                             
                tmr_registers(1)(730)    <= not(global_tmr_voter(1)(729));                                                             
                tmr_registers(2)(730)    <= not(global_tmr_voter(2)(729));                                                             
 
                tmr_registers(0)(731)    <= not(global_tmr_voter(0)(730));                                                             
                tmr_registers(1)(731)    <= not(global_tmr_voter(1)(730));                                                             
                tmr_registers(2)(731)    <= not(global_tmr_voter(2)(730));                                                             
 
                tmr_registers(0)(732)    <= not(global_tmr_voter(0)(731));                                                             
                tmr_registers(1)(732)    <= not(global_tmr_voter(1)(731));                                                             
                tmr_registers(2)(732)    <= not(global_tmr_voter(2)(731));                                                             
 
                tmr_registers(0)(733)    <= not(global_tmr_voter(0)(732));                                                             
                tmr_registers(1)(733)    <= not(global_tmr_voter(1)(732));                                                             
                tmr_registers(2)(733)    <= not(global_tmr_voter(2)(732));                                                             
 
                tmr_registers(0)(734)    <= not(global_tmr_voter(0)(733));                                                             
                tmr_registers(1)(734)    <= not(global_tmr_voter(1)(733));                                                             
                tmr_registers(2)(734)    <= not(global_tmr_voter(2)(733));                                                             
 
                tmr_registers(0)(735)    <= not(global_tmr_voter(0)(734));                                                             
                tmr_registers(1)(735)    <= not(global_tmr_voter(1)(734));                                                             
                tmr_registers(2)(735)    <= not(global_tmr_voter(2)(734));                                                             
 
                tmr_registers(0)(736)    <= not(global_tmr_voter(0)(735));                                                             
                tmr_registers(1)(736)    <= not(global_tmr_voter(1)(735));                                                             
                tmr_registers(2)(736)    <= not(global_tmr_voter(2)(735));                                                             
 
                tmr_registers(0)(737)    <= not(global_tmr_voter(0)(736));                                                             
                tmr_registers(1)(737)    <= not(global_tmr_voter(1)(736));                                                             
                tmr_registers(2)(737)    <= not(global_tmr_voter(2)(736));                                                             
 
                tmr_registers(0)(738)    <= not(global_tmr_voter(0)(737));                                                             
                tmr_registers(1)(738)    <= not(global_tmr_voter(1)(737));                                                             
                tmr_registers(2)(738)    <= not(global_tmr_voter(2)(737));                                                             
 
                tmr_registers(0)(739)    <= not(global_tmr_voter(0)(738));                                                             
                tmr_registers(1)(739)    <= not(global_tmr_voter(1)(738));                                                             
                tmr_registers(2)(739)    <= not(global_tmr_voter(2)(738));                                                             
 
                tmr_registers(0)(740)    <= not(global_tmr_voter(0)(739));                                                             
                tmr_registers(1)(740)    <= not(global_tmr_voter(1)(739));                                                             
                tmr_registers(2)(740)    <= not(global_tmr_voter(2)(739));                                                             
 
                tmr_registers(0)(741)    <= not(global_tmr_voter(0)(740));                                                             
                tmr_registers(1)(741)    <= not(global_tmr_voter(1)(740));                                                             
                tmr_registers(2)(741)    <= not(global_tmr_voter(2)(740));                                                             
 
                tmr_registers(0)(742)    <= not(global_tmr_voter(0)(741));                                                             
                tmr_registers(1)(742)    <= not(global_tmr_voter(1)(741));                                                             
                tmr_registers(2)(742)    <= not(global_tmr_voter(2)(741));                                                             
 
                tmr_registers(0)(743)    <= not(global_tmr_voter(0)(742));                                                             
                tmr_registers(1)(743)    <= not(global_tmr_voter(1)(742));                                                             
                tmr_registers(2)(743)    <= not(global_tmr_voter(2)(742));                                                             
 
                tmr_registers(0)(744)    <= not(global_tmr_voter(0)(743));                                                             
                tmr_registers(1)(744)    <= not(global_tmr_voter(1)(743));                                                             
                tmr_registers(2)(744)    <= not(global_tmr_voter(2)(743));                                                             
 
                tmr_registers(0)(745)    <= not(global_tmr_voter(0)(744));                                                             
                tmr_registers(1)(745)    <= not(global_tmr_voter(1)(744));                                                             
                tmr_registers(2)(745)    <= not(global_tmr_voter(2)(744));                                                             
 
                tmr_registers(0)(746)    <= not(global_tmr_voter(0)(745));                                                             
                tmr_registers(1)(746)    <= not(global_tmr_voter(1)(745));                                                             
                tmr_registers(2)(746)    <= not(global_tmr_voter(2)(745));                                                             
 
                tmr_registers(0)(747)    <= not(global_tmr_voter(0)(746));                                                             
                tmr_registers(1)(747)    <= not(global_tmr_voter(1)(746));                                                             
                tmr_registers(2)(747)    <= not(global_tmr_voter(2)(746));                                                             
 
                tmr_registers(0)(748)    <= not(global_tmr_voter(0)(747));                                                             
                tmr_registers(1)(748)    <= not(global_tmr_voter(1)(747));                                                             
                tmr_registers(2)(748)    <= not(global_tmr_voter(2)(747));                                                             
 
                tmr_registers(0)(749)    <= not(global_tmr_voter(0)(748));                                                             
                tmr_registers(1)(749)    <= not(global_tmr_voter(1)(748));                                                             
                tmr_registers(2)(749)    <= not(global_tmr_voter(2)(748));                                                             
 
                tmr_registers(0)(750)    <= not(global_tmr_voter(0)(749));                                                             
                tmr_registers(1)(750)    <= not(global_tmr_voter(1)(749));                                                             
                tmr_registers(2)(750)    <= not(global_tmr_voter(2)(749));                                                             
 
                tmr_registers(0)(751)    <= not(global_tmr_voter(0)(750));                                                             
                tmr_registers(1)(751)    <= not(global_tmr_voter(1)(750));                                                             
                tmr_registers(2)(751)    <= not(global_tmr_voter(2)(750));                                                             
 
                tmr_registers(0)(752)    <= not(global_tmr_voter(0)(751));                                                             
                tmr_registers(1)(752)    <= not(global_tmr_voter(1)(751));                                                             
                tmr_registers(2)(752)    <= not(global_tmr_voter(2)(751));                                                             
 
                tmr_registers(0)(753)    <= not(global_tmr_voter(0)(752));                                                             
                tmr_registers(1)(753)    <= not(global_tmr_voter(1)(752));                                                             
                tmr_registers(2)(753)    <= not(global_tmr_voter(2)(752));                                                             
 
                tmr_registers(0)(754)    <= not(global_tmr_voter(0)(753));                                                             
                tmr_registers(1)(754)    <= not(global_tmr_voter(1)(753));                                                             
                tmr_registers(2)(754)    <= not(global_tmr_voter(2)(753));                                                             
 
                tmr_registers(0)(755)    <= not(global_tmr_voter(0)(754));                                                             
                tmr_registers(1)(755)    <= not(global_tmr_voter(1)(754));                                                             
                tmr_registers(2)(755)    <= not(global_tmr_voter(2)(754));                                                             
 
                tmr_registers(0)(756)    <= not(global_tmr_voter(0)(755));                                                             
                tmr_registers(1)(756)    <= not(global_tmr_voter(1)(755));                                                             
                tmr_registers(2)(756)    <= not(global_tmr_voter(2)(755));                                                             
 
                tmr_registers(0)(757)    <= not(global_tmr_voter(0)(756));                                                             
                tmr_registers(1)(757)    <= not(global_tmr_voter(1)(756));                                                             
                tmr_registers(2)(757)    <= not(global_tmr_voter(2)(756));                                                             
 
                tmr_registers(0)(758)    <= not(global_tmr_voter(0)(757));                                                             
                tmr_registers(1)(758)    <= not(global_tmr_voter(1)(757));                                                             
                tmr_registers(2)(758)    <= not(global_tmr_voter(2)(757));                                                             
 
                tmr_registers(0)(759)    <= not(global_tmr_voter(0)(758));                                                             
                tmr_registers(1)(759)    <= not(global_tmr_voter(1)(758));                                                             
                tmr_registers(2)(759)    <= not(global_tmr_voter(2)(758));                                                             
 
                tmr_registers(0)(760)    <= not(global_tmr_voter(0)(759));                                                             
                tmr_registers(1)(760)    <= not(global_tmr_voter(1)(759));                                                             
                tmr_registers(2)(760)    <= not(global_tmr_voter(2)(759));                                                             
 
                tmr_registers(0)(761)    <= not(global_tmr_voter(0)(760));                                                             
                tmr_registers(1)(761)    <= not(global_tmr_voter(1)(760));                                                             
                tmr_registers(2)(761)    <= not(global_tmr_voter(2)(760));                                                             
 
                tmr_registers(0)(762)    <= not(global_tmr_voter(0)(761));                                                             
                tmr_registers(1)(762)    <= not(global_tmr_voter(1)(761));                                                             
                tmr_registers(2)(762)    <= not(global_tmr_voter(2)(761));                                                             
 
                tmr_registers(0)(763)    <= not(global_tmr_voter(0)(762));                                                             
                tmr_registers(1)(763)    <= not(global_tmr_voter(1)(762));                                                             
                tmr_registers(2)(763)    <= not(global_tmr_voter(2)(762));                                                             
 
                tmr_registers(0)(764)    <= not(global_tmr_voter(0)(763));                                                             
                tmr_registers(1)(764)    <= not(global_tmr_voter(1)(763));                                                             
                tmr_registers(2)(764)    <= not(global_tmr_voter(2)(763));                                                             
 
                tmr_registers(0)(765)    <= not(global_tmr_voter(0)(764));                                                             
                tmr_registers(1)(765)    <= not(global_tmr_voter(1)(764));                                                             
                tmr_registers(2)(765)    <= not(global_tmr_voter(2)(764));                                                             
 
                tmr_registers(0)(766)    <= not(global_tmr_voter(0)(765));                                                             
                tmr_registers(1)(766)    <= not(global_tmr_voter(1)(765));                                                             
                tmr_registers(2)(766)    <= not(global_tmr_voter(2)(765));                                                             
 
                tmr_registers(0)(767)    <= not(global_tmr_voter(0)(766));                                                             
                tmr_registers(1)(767)    <= not(global_tmr_voter(1)(766));                                                             
                tmr_registers(2)(767)    <= not(global_tmr_voter(2)(766));                                                             
 
                tmr_registers(0)(768)    <= not(global_tmr_voter(0)(767));                                                             
                tmr_registers(1)(768)    <= not(global_tmr_voter(1)(767));                                                             
                tmr_registers(2)(768)    <= not(global_tmr_voter(2)(767));                                                             
 
                tmr_registers(0)(769)    <= not(global_tmr_voter(0)(768));                                                             
                tmr_registers(1)(769)    <= not(global_tmr_voter(1)(768));                                                             
                tmr_registers(2)(769)    <= not(global_tmr_voter(2)(768));                                                             
 
                tmr_registers(0)(770)    <= not(global_tmr_voter(0)(769));                                                             
                tmr_registers(1)(770)    <= not(global_tmr_voter(1)(769));                                                             
                tmr_registers(2)(770)    <= not(global_tmr_voter(2)(769));                                                             
 
                tmr_registers(0)(771)    <= not(global_tmr_voter(0)(770));                                                             
                tmr_registers(1)(771)    <= not(global_tmr_voter(1)(770));                                                             
                tmr_registers(2)(771)    <= not(global_tmr_voter(2)(770));                                                             
 
                tmr_registers(0)(772)    <= not(global_tmr_voter(0)(771));                                                             
                tmr_registers(1)(772)    <= not(global_tmr_voter(1)(771));                                                             
                tmr_registers(2)(772)    <= not(global_tmr_voter(2)(771));                                                             
 
                tmr_registers(0)(773)    <= not(global_tmr_voter(0)(772));                                                             
                tmr_registers(1)(773)    <= not(global_tmr_voter(1)(772));                                                             
                tmr_registers(2)(773)    <= not(global_tmr_voter(2)(772));                                                             
 
                tmr_registers(0)(774)    <= not(global_tmr_voter(0)(773));                                                             
                tmr_registers(1)(774)    <= not(global_tmr_voter(1)(773));                                                             
                tmr_registers(2)(774)    <= not(global_tmr_voter(2)(773));                                                             
 
                tmr_registers(0)(775)    <= not(global_tmr_voter(0)(774));                                                             
                tmr_registers(1)(775)    <= not(global_tmr_voter(1)(774));                                                             
                tmr_registers(2)(775)    <= not(global_tmr_voter(2)(774));                                                             
 
                tmr_registers(0)(776)    <= not(global_tmr_voter(0)(775));                                                             
                tmr_registers(1)(776)    <= not(global_tmr_voter(1)(775));                                                             
                tmr_registers(2)(776)    <= not(global_tmr_voter(2)(775));                                                             
 
                tmr_registers(0)(777)    <= not(global_tmr_voter(0)(776));                                                             
                tmr_registers(1)(777)    <= not(global_tmr_voter(1)(776));                                                             
                tmr_registers(2)(777)    <= not(global_tmr_voter(2)(776));                                                             
 
                tmr_registers(0)(778)    <= not(global_tmr_voter(0)(777));                                                             
                tmr_registers(1)(778)    <= not(global_tmr_voter(1)(777));                                                             
                tmr_registers(2)(778)    <= not(global_tmr_voter(2)(777));                                                             
 
                tmr_registers(0)(779)    <= not(global_tmr_voter(0)(778));                                                             
                tmr_registers(1)(779)    <= not(global_tmr_voter(1)(778));                                                             
                tmr_registers(2)(779)    <= not(global_tmr_voter(2)(778));                                                             
 
                tmr_registers(0)(780)    <= not(global_tmr_voter(0)(779));                                                             
                tmr_registers(1)(780)    <= not(global_tmr_voter(1)(779));                                                             
                tmr_registers(2)(780)    <= not(global_tmr_voter(2)(779));                                                             
 
                tmr_registers(0)(781)    <= not(global_tmr_voter(0)(780));                                                             
                tmr_registers(1)(781)    <= not(global_tmr_voter(1)(780));                                                             
                tmr_registers(2)(781)    <= not(global_tmr_voter(2)(780));                                                             
 
                tmr_registers(0)(782)    <= not(global_tmr_voter(0)(781));                                                             
                tmr_registers(1)(782)    <= not(global_tmr_voter(1)(781));                                                             
                tmr_registers(2)(782)    <= not(global_tmr_voter(2)(781));                                                             
 
                tmr_registers(0)(783)    <= not(global_tmr_voter(0)(782));                                                             
                tmr_registers(1)(783)    <= not(global_tmr_voter(1)(782));                                                             
                tmr_registers(2)(783)    <= not(global_tmr_voter(2)(782));                                                             
 
                tmr_registers(0)(784)    <= not(global_tmr_voter(0)(783));                                                             
                tmr_registers(1)(784)    <= not(global_tmr_voter(1)(783));                                                             
                tmr_registers(2)(784)    <= not(global_tmr_voter(2)(783));                                                             
 
                tmr_registers(0)(785)    <= not(global_tmr_voter(0)(784));                                                             
                tmr_registers(1)(785)    <= not(global_tmr_voter(1)(784));                                                             
                tmr_registers(2)(785)    <= not(global_tmr_voter(2)(784));                                                             
 
                tmr_registers(0)(786)    <= not(global_tmr_voter(0)(785));                                                             
                tmr_registers(1)(786)    <= not(global_tmr_voter(1)(785));                                                             
                tmr_registers(2)(786)    <= not(global_tmr_voter(2)(785));                                                             
 
                tmr_registers(0)(787)    <= not(global_tmr_voter(0)(786));                                                             
                tmr_registers(1)(787)    <= not(global_tmr_voter(1)(786));                                                             
                tmr_registers(2)(787)    <= not(global_tmr_voter(2)(786));                                                             
 
                tmr_registers(0)(788)    <= not(global_tmr_voter(0)(787));                                                             
                tmr_registers(1)(788)    <= not(global_tmr_voter(1)(787));                                                             
                tmr_registers(2)(788)    <= not(global_tmr_voter(2)(787));                                                             
 
                tmr_registers(0)(789)    <= not(global_tmr_voter(0)(788));                                                             
                tmr_registers(1)(789)    <= not(global_tmr_voter(1)(788));                                                             
                tmr_registers(2)(789)    <= not(global_tmr_voter(2)(788));                                                             
 
                tmr_registers(0)(790)    <= not(global_tmr_voter(0)(789));                                                             
                tmr_registers(1)(790)    <= not(global_tmr_voter(1)(789));                                                             
                tmr_registers(2)(790)    <= not(global_tmr_voter(2)(789));                                                             
 
                tmr_registers(0)(791)    <= not(global_tmr_voter(0)(790));                                                             
                tmr_registers(1)(791)    <= not(global_tmr_voter(1)(790));                                                             
                tmr_registers(2)(791)    <= not(global_tmr_voter(2)(790));                                                             
 
                tmr_registers(0)(792)    <= not(global_tmr_voter(0)(791));                                                             
                tmr_registers(1)(792)    <= not(global_tmr_voter(1)(791));                                                             
                tmr_registers(2)(792)    <= not(global_tmr_voter(2)(791));                                                             
 
                tmr_registers(0)(793)    <= not(global_tmr_voter(0)(792));                                                             
                tmr_registers(1)(793)    <= not(global_tmr_voter(1)(792));                                                             
                tmr_registers(2)(793)    <= not(global_tmr_voter(2)(792));                                                             
 
                tmr_registers(0)(794)    <= not(global_tmr_voter(0)(793));                                                             
                tmr_registers(1)(794)    <= not(global_tmr_voter(1)(793));                                                             
                tmr_registers(2)(794)    <= not(global_tmr_voter(2)(793));                                                             
 
                tmr_registers(0)(795)    <= not(global_tmr_voter(0)(794));                                                             
                tmr_registers(1)(795)    <= not(global_tmr_voter(1)(794));                                                             
                tmr_registers(2)(795)    <= not(global_tmr_voter(2)(794));                                                             
 
                tmr_registers(0)(796)    <= not(global_tmr_voter(0)(795));                                                             
                tmr_registers(1)(796)    <= not(global_tmr_voter(1)(795));                                                             
                tmr_registers(2)(796)    <= not(global_tmr_voter(2)(795));                                                             
 
                tmr_registers(0)(797)    <= not(global_tmr_voter(0)(796));                                                             
                tmr_registers(1)(797)    <= not(global_tmr_voter(1)(796));                                                             
                tmr_registers(2)(797)    <= not(global_tmr_voter(2)(796));                                                             
 
                tmr_registers(0)(798)    <= not(global_tmr_voter(0)(797));                                                             
                tmr_registers(1)(798)    <= not(global_tmr_voter(1)(797));                                                             
                tmr_registers(2)(798)    <= not(global_tmr_voter(2)(797));                                                             
 
                tmr_registers(0)(799)    <= not(global_tmr_voter(0)(798));                                                             
                tmr_registers(1)(799)    <= not(global_tmr_voter(1)(798));                                                             
                tmr_registers(2)(799)    <= not(global_tmr_voter(2)(798));                                                             
 
                tmr_registers(0)(800)    <= not(global_tmr_voter(0)(799));                                                             
                tmr_registers(1)(800)    <= not(global_tmr_voter(1)(799));                                                             
                tmr_registers(2)(800)    <= not(global_tmr_voter(2)(799));                                                             
 
                tmr_registers(0)(801)    <= not(global_tmr_voter(0)(800));                                                             
                tmr_registers(1)(801)    <= not(global_tmr_voter(1)(800));                                                             
                tmr_registers(2)(801)    <= not(global_tmr_voter(2)(800));                                                             
 
                tmr_registers(0)(802)    <= not(global_tmr_voter(0)(801));                                                             
                tmr_registers(1)(802)    <= not(global_tmr_voter(1)(801));                                                             
                tmr_registers(2)(802)    <= not(global_tmr_voter(2)(801));                                                             
 
                tmr_registers(0)(803)    <= not(global_tmr_voter(0)(802));                                                             
                tmr_registers(1)(803)    <= not(global_tmr_voter(1)(802));                                                             
                tmr_registers(2)(803)    <= not(global_tmr_voter(2)(802));                                                             
 
                tmr_registers(0)(804)    <= not(global_tmr_voter(0)(803));                                                             
                tmr_registers(1)(804)    <= not(global_tmr_voter(1)(803));                                                             
                tmr_registers(2)(804)    <= not(global_tmr_voter(2)(803));                                                             
 
                tmr_registers(0)(805)    <= not(global_tmr_voter(0)(804));                                                             
                tmr_registers(1)(805)    <= not(global_tmr_voter(1)(804));                                                             
                tmr_registers(2)(805)    <= not(global_tmr_voter(2)(804));                                                             
 
                tmr_registers(0)(806)    <= not(global_tmr_voter(0)(805));                                                             
                tmr_registers(1)(806)    <= not(global_tmr_voter(1)(805));                                                             
                tmr_registers(2)(806)    <= not(global_tmr_voter(2)(805));                                                             
 
                tmr_registers(0)(807)    <= not(global_tmr_voter(0)(806));                                                             
                tmr_registers(1)(807)    <= not(global_tmr_voter(1)(806));                                                             
                tmr_registers(2)(807)    <= not(global_tmr_voter(2)(806));                                                             
 
                tmr_registers(0)(808)    <= not(global_tmr_voter(0)(807));                                                             
                tmr_registers(1)(808)    <= not(global_tmr_voter(1)(807));                                                             
                tmr_registers(2)(808)    <= not(global_tmr_voter(2)(807));                                                             
 
                tmr_registers(0)(809)    <= not(global_tmr_voter(0)(808));                                                             
                tmr_registers(1)(809)    <= not(global_tmr_voter(1)(808));                                                             
                tmr_registers(2)(809)    <= not(global_tmr_voter(2)(808));                                                             
 
                tmr_registers(0)(810)    <= not(global_tmr_voter(0)(809));                                                             
                tmr_registers(1)(810)    <= not(global_tmr_voter(1)(809));                                                             
                tmr_registers(2)(810)    <= not(global_tmr_voter(2)(809));                                                             
 
                tmr_registers(0)(811)    <= not(global_tmr_voter(0)(810));                                                             
                tmr_registers(1)(811)    <= not(global_tmr_voter(1)(810));                                                             
                tmr_registers(2)(811)    <= not(global_tmr_voter(2)(810));                                                             
 
                tmr_registers(0)(812)    <= not(global_tmr_voter(0)(811));                                                             
                tmr_registers(1)(812)    <= not(global_tmr_voter(1)(811));                                                             
                tmr_registers(2)(812)    <= not(global_tmr_voter(2)(811));                                                             
 
                tmr_registers(0)(813)    <= not(global_tmr_voter(0)(812));                                                             
                tmr_registers(1)(813)    <= not(global_tmr_voter(1)(812));                                                             
                tmr_registers(2)(813)    <= not(global_tmr_voter(2)(812));                                                             
 
                tmr_registers(0)(814)    <= not(global_tmr_voter(0)(813));                                                             
                tmr_registers(1)(814)    <= not(global_tmr_voter(1)(813));                                                             
                tmr_registers(2)(814)    <= not(global_tmr_voter(2)(813));                                                             
 
                tmr_registers(0)(815)    <= not(global_tmr_voter(0)(814));                                                             
                tmr_registers(1)(815)    <= not(global_tmr_voter(1)(814));                                                             
                tmr_registers(2)(815)    <= not(global_tmr_voter(2)(814));                                                             
 
                tmr_registers(0)(816)    <= not(global_tmr_voter(0)(815));                                                             
                tmr_registers(1)(816)    <= not(global_tmr_voter(1)(815));                                                             
                tmr_registers(2)(816)    <= not(global_tmr_voter(2)(815));                                                             
 
                tmr_registers(0)(817)    <= not(global_tmr_voter(0)(816));                                                             
                tmr_registers(1)(817)    <= not(global_tmr_voter(1)(816));                                                             
                tmr_registers(2)(817)    <= not(global_tmr_voter(2)(816));                                                             
 
                tmr_registers(0)(818)    <= not(global_tmr_voter(0)(817));                                                             
                tmr_registers(1)(818)    <= not(global_tmr_voter(1)(817));                                                             
                tmr_registers(2)(818)    <= not(global_tmr_voter(2)(817));                                                             
 
                tmr_registers(0)(819)    <= not(global_tmr_voter(0)(818));                                                             
                tmr_registers(1)(819)    <= not(global_tmr_voter(1)(818));                                                             
                tmr_registers(2)(819)    <= not(global_tmr_voter(2)(818));                                                             
 
                tmr_registers(0)(820)    <= not(global_tmr_voter(0)(819));                                                             
                tmr_registers(1)(820)    <= not(global_tmr_voter(1)(819));                                                             
                tmr_registers(2)(820)    <= not(global_tmr_voter(2)(819));                                                             
 
                tmr_registers(0)(821)    <= not(global_tmr_voter(0)(820));                                                             
                tmr_registers(1)(821)    <= not(global_tmr_voter(1)(820));                                                             
                tmr_registers(2)(821)    <= not(global_tmr_voter(2)(820));                                                             
 
                tmr_registers(0)(822)    <= not(global_tmr_voter(0)(821));                                                             
                tmr_registers(1)(822)    <= not(global_tmr_voter(1)(821));                                                             
                tmr_registers(2)(822)    <= not(global_tmr_voter(2)(821));                                                             
 
                tmr_registers(0)(823)    <= not(global_tmr_voter(0)(822));                                                             
                tmr_registers(1)(823)    <= not(global_tmr_voter(1)(822));                                                             
                tmr_registers(2)(823)    <= not(global_tmr_voter(2)(822));                                                             
 
                tmr_registers(0)(824)    <= not(global_tmr_voter(0)(823));                                                             
                tmr_registers(1)(824)    <= not(global_tmr_voter(1)(823));                                                             
                tmr_registers(2)(824)    <= not(global_tmr_voter(2)(823));                                                             
 
                tmr_registers(0)(825)    <= not(global_tmr_voter(0)(824));                                                             
                tmr_registers(1)(825)    <= not(global_tmr_voter(1)(824));                                                             
                tmr_registers(2)(825)    <= not(global_tmr_voter(2)(824));                                                             
 
                tmr_registers(0)(826)    <= not(global_tmr_voter(0)(825));                                                             
                tmr_registers(1)(826)    <= not(global_tmr_voter(1)(825));                                                             
                tmr_registers(2)(826)    <= not(global_tmr_voter(2)(825));                                                             
 
                tmr_registers(0)(827)    <= not(global_tmr_voter(0)(826));                                                             
                tmr_registers(1)(827)    <= not(global_tmr_voter(1)(826));                                                             
                tmr_registers(2)(827)    <= not(global_tmr_voter(2)(826));                                                             
 
                tmr_registers(0)(828)    <= not(global_tmr_voter(0)(827));                                                             
                tmr_registers(1)(828)    <= not(global_tmr_voter(1)(827));                                                             
                tmr_registers(2)(828)    <= not(global_tmr_voter(2)(827));                                                             
 
                tmr_registers(0)(829)    <= not(global_tmr_voter(0)(828));                                                             
                tmr_registers(1)(829)    <= not(global_tmr_voter(1)(828));                                                             
                tmr_registers(2)(829)    <= not(global_tmr_voter(2)(828));                                                             
 
                tmr_registers(0)(830)    <= not(global_tmr_voter(0)(829));                                                             
                tmr_registers(1)(830)    <= not(global_tmr_voter(1)(829));                                                             
                tmr_registers(2)(830)    <= not(global_tmr_voter(2)(829));                                                             
 
                tmr_registers(0)(831)    <= not(global_tmr_voter(0)(830));                                                             
                tmr_registers(1)(831)    <= not(global_tmr_voter(1)(830));                                                             
                tmr_registers(2)(831)    <= not(global_tmr_voter(2)(830));                                                             
 
                tmr_registers(0)(832)    <= not(global_tmr_voter(0)(831));                                                             
                tmr_registers(1)(832)    <= not(global_tmr_voter(1)(831));                                                             
                tmr_registers(2)(832)    <= not(global_tmr_voter(2)(831));                                                             
 
                tmr_registers(0)(833)    <= not(global_tmr_voter(0)(832));                                                             
                tmr_registers(1)(833)    <= not(global_tmr_voter(1)(832));                                                             
                tmr_registers(2)(833)    <= not(global_tmr_voter(2)(832));                                                             
 
                tmr_registers(0)(834)    <= not(global_tmr_voter(0)(833));                                                             
                tmr_registers(1)(834)    <= not(global_tmr_voter(1)(833));                                                             
                tmr_registers(2)(834)    <= not(global_tmr_voter(2)(833));                                                             
 
                tmr_registers(0)(835)    <= not(global_tmr_voter(0)(834));                                                             
                tmr_registers(1)(835)    <= not(global_tmr_voter(1)(834));                                                             
                tmr_registers(2)(835)    <= not(global_tmr_voter(2)(834));                                                             
 
                tmr_registers(0)(836)    <= not(global_tmr_voter(0)(835));                                                             
                tmr_registers(1)(836)    <= not(global_tmr_voter(1)(835));                                                             
                tmr_registers(2)(836)    <= not(global_tmr_voter(2)(835));                                                             
 
                tmr_registers(0)(837)    <= not(global_tmr_voter(0)(836));                                                             
                tmr_registers(1)(837)    <= not(global_tmr_voter(1)(836));                                                             
                tmr_registers(2)(837)    <= not(global_tmr_voter(2)(836));                                                             
 
                tmr_registers(0)(838)    <= not(global_tmr_voter(0)(837));                                                             
                tmr_registers(1)(838)    <= not(global_tmr_voter(1)(837));                                                             
                tmr_registers(2)(838)    <= not(global_tmr_voter(2)(837));                                                             
 
                tmr_registers(0)(839)    <= not(global_tmr_voter(0)(838));                                                             
                tmr_registers(1)(839)    <= not(global_tmr_voter(1)(838));                                                             
                tmr_registers(2)(839)    <= not(global_tmr_voter(2)(838));                                                             
 
                tmr_registers(0)(840)    <= not(global_tmr_voter(0)(839));                                                             
                tmr_registers(1)(840)    <= not(global_tmr_voter(1)(839));                                                             
                tmr_registers(2)(840)    <= not(global_tmr_voter(2)(839));                                                             
 
                tmr_registers(0)(841)    <= not(global_tmr_voter(0)(840));                                                             
                tmr_registers(1)(841)    <= not(global_tmr_voter(1)(840));                                                             
                tmr_registers(2)(841)    <= not(global_tmr_voter(2)(840));                                                             
 
                tmr_registers(0)(842)    <= not(global_tmr_voter(0)(841));                                                             
                tmr_registers(1)(842)    <= not(global_tmr_voter(1)(841));                                                             
                tmr_registers(2)(842)    <= not(global_tmr_voter(2)(841));                                                             
 
                tmr_registers(0)(843)    <= not(global_tmr_voter(0)(842));                                                             
                tmr_registers(1)(843)    <= not(global_tmr_voter(1)(842));                                                             
                tmr_registers(2)(843)    <= not(global_tmr_voter(2)(842));                                                             
 
                tmr_registers(0)(844)    <= not(global_tmr_voter(0)(843));                                                             
                tmr_registers(1)(844)    <= not(global_tmr_voter(1)(843));                                                             
                tmr_registers(2)(844)    <= not(global_tmr_voter(2)(843));                                                             
 
                tmr_registers(0)(845)    <= not(global_tmr_voter(0)(844));                                                             
                tmr_registers(1)(845)    <= not(global_tmr_voter(1)(844));                                                             
                tmr_registers(2)(845)    <= not(global_tmr_voter(2)(844));                                                             
 
                tmr_registers(0)(846)    <= not(global_tmr_voter(0)(845));                                                             
                tmr_registers(1)(846)    <= not(global_tmr_voter(1)(845));                                                             
                tmr_registers(2)(846)    <= not(global_tmr_voter(2)(845));                                                             
 
                tmr_registers(0)(847)    <= not(global_tmr_voter(0)(846));                                                             
                tmr_registers(1)(847)    <= not(global_tmr_voter(1)(846));                                                             
                tmr_registers(2)(847)    <= not(global_tmr_voter(2)(846));                                                             
 
                tmr_registers(0)(848)    <= not(global_tmr_voter(0)(847));                                                             
                tmr_registers(1)(848)    <= not(global_tmr_voter(1)(847));                                                             
                tmr_registers(2)(848)    <= not(global_tmr_voter(2)(847));                                                             
 
                tmr_registers(0)(849)    <= not(global_tmr_voter(0)(848));                                                             
                tmr_registers(1)(849)    <= not(global_tmr_voter(1)(848));                                                             
                tmr_registers(2)(849)    <= not(global_tmr_voter(2)(848));                                                             
 
                tmr_registers(0)(850)    <= not(global_tmr_voter(0)(849));                                                             
                tmr_registers(1)(850)    <= not(global_tmr_voter(1)(849));                                                             
                tmr_registers(2)(850)    <= not(global_tmr_voter(2)(849));                                                             
 
                tmr_registers(0)(851)    <= not(global_tmr_voter(0)(850));                                                             
                tmr_registers(1)(851)    <= not(global_tmr_voter(1)(850));                                                             
                tmr_registers(2)(851)    <= not(global_tmr_voter(2)(850));                                                             
 
                tmr_registers(0)(852)    <= not(global_tmr_voter(0)(851));                                                             
                tmr_registers(1)(852)    <= not(global_tmr_voter(1)(851));                                                             
                tmr_registers(2)(852)    <= not(global_tmr_voter(2)(851));                                                             
 
                tmr_registers(0)(853)    <= not(global_tmr_voter(0)(852));                                                             
                tmr_registers(1)(853)    <= not(global_tmr_voter(1)(852));                                                             
                tmr_registers(2)(853)    <= not(global_tmr_voter(2)(852));                                                             
 
                tmr_registers(0)(854)    <= not(global_tmr_voter(0)(853));                                                             
                tmr_registers(1)(854)    <= not(global_tmr_voter(1)(853));                                                             
                tmr_registers(2)(854)    <= not(global_tmr_voter(2)(853));                                                             
 
                tmr_registers(0)(855)    <= not(global_tmr_voter(0)(854));                                                             
                tmr_registers(1)(855)    <= not(global_tmr_voter(1)(854));                                                             
                tmr_registers(2)(855)    <= not(global_tmr_voter(2)(854));                                                             
 
                tmr_registers(0)(856)    <= not(global_tmr_voter(0)(855));                                                             
                tmr_registers(1)(856)    <= not(global_tmr_voter(1)(855));                                                             
                tmr_registers(2)(856)    <= not(global_tmr_voter(2)(855));                                                             
 
                tmr_registers(0)(857)    <= not(global_tmr_voter(0)(856));                                                             
                tmr_registers(1)(857)    <= not(global_tmr_voter(1)(856));                                                             
                tmr_registers(2)(857)    <= not(global_tmr_voter(2)(856));                                                             
 
                tmr_registers(0)(858)    <= not(global_tmr_voter(0)(857));                                                             
                tmr_registers(1)(858)    <= not(global_tmr_voter(1)(857));                                                             
                tmr_registers(2)(858)    <= not(global_tmr_voter(2)(857));                                                             
 
                tmr_registers(0)(859)    <= not(global_tmr_voter(0)(858));                                                             
                tmr_registers(1)(859)    <= not(global_tmr_voter(1)(858));                                                             
                tmr_registers(2)(859)    <= not(global_tmr_voter(2)(858));                                                             
 
                tmr_registers(0)(860)    <= not(global_tmr_voter(0)(859));                                                             
                tmr_registers(1)(860)    <= not(global_tmr_voter(1)(859));                                                             
                tmr_registers(2)(860)    <= not(global_tmr_voter(2)(859));                                                             
 
                tmr_registers(0)(861)    <= not(global_tmr_voter(0)(860));                                                             
                tmr_registers(1)(861)    <= not(global_tmr_voter(1)(860));                                                             
                tmr_registers(2)(861)    <= not(global_tmr_voter(2)(860));                                                             
 
                tmr_registers(0)(862)    <= not(global_tmr_voter(0)(861));                                                             
                tmr_registers(1)(862)    <= not(global_tmr_voter(1)(861));                                                             
                tmr_registers(2)(862)    <= not(global_tmr_voter(2)(861));                                                             
 
                tmr_registers(0)(863)    <= not(global_tmr_voter(0)(862));                                                             
                tmr_registers(1)(863)    <= not(global_tmr_voter(1)(862));                                                             
                tmr_registers(2)(863)    <= not(global_tmr_voter(2)(862));                                                             
 
                tmr_registers(0)(864)    <= not(global_tmr_voter(0)(863));                                                             
                tmr_registers(1)(864)    <= not(global_tmr_voter(1)(863));                                                             
                tmr_registers(2)(864)    <= not(global_tmr_voter(2)(863));                                                             
 
                tmr_registers(0)(865)    <= not(global_tmr_voter(0)(864));                                                             
                tmr_registers(1)(865)    <= not(global_tmr_voter(1)(864));                                                             
                tmr_registers(2)(865)    <= not(global_tmr_voter(2)(864));                                                             
 
                tmr_registers(0)(866)    <= not(global_tmr_voter(0)(865));                                                             
                tmr_registers(1)(866)    <= not(global_tmr_voter(1)(865));                                                             
                tmr_registers(2)(866)    <= not(global_tmr_voter(2)(865));                                                             
 
                tmr_registers(0)(867)    <= not(global_tmr_voter(0)(866));                                                             
                tmr_registers(1)(867)    <= not(global_tmr_voter(1)(866));                                                             
                tmr_registers(2)(867)    <= not(global_tmr_voter(2)(866));                                                             
 
                tmr_registers(0)(868)    <= not(global_tmr_voter(0)(867));                                                             
                tmr_registers(1)(868)    <= not(global_tmr_voter(1)(867));                                                             
                tmr_registers(2)(868)    <= not(global_tmr_voter(2)(867));                                                             
 
                tmr_registers(0)(869)    <= not(global_tmr_voter(0)(868));                                                             
                tmr_registers(1)(869)    <= not(global_tmr_voter(1)(868));                                                             
                tmr_registers(2)(869)    <= not(global_tmr_voter(2)(868));                                                             
 
                tmr_registers(0)(870)    <= not(global_tmr_voter(0)(869));                                                             
                tmr_registers(1)(870)    <= not(global_tmr_voter(1)(869));                                                             
                tmr_registers(2)(870)    <= not(global_tmr_voter(2)(869));                                                             
 
                tmr_registers(0)(871)    <= not(global_tmr_voter(0)(870));                                                             
                tmr_registers(1)(871)    <= not(global_tmr_voter(1)(870));                                                             
                tmr_registers(2)(871)    <= not(global_tmr_voter(2)(870));                                                             
 
                tmr_registers(0)(872)    <= not(global_tmr_voter(0)(871));                                                             
                tmr_registers(1)(872)    <= not(global_tmr_voter(1)(871));                                                             
                tmr_registers(2)(872)    <= not(global_tmr_voter(2)(871));                                                             
 
                tmr_registers(0)(873)    <= not(global_tmr_voter(0)(872));                                                             
                tmr_registers(1)(873)    <= not(global_tmr_voter(1)(872));                                                             
                tmr_registers(2)(873)    <= not(global_tmr_voter(2)(872));                                                             
 
                tmr_registers(0)(874)    <= not(global_tmr_voter(0)(873));                                                             
                tmr_registers(1)(874)    <= not(global_tmr_voter(1)(873));                                                             
                tmr_registers(2)(874)    <= not(global_tmr_voter(2)(873));                                                             
 
                tmr_registers(0)(875)    <= not(global_tmr_voter(0)(874));                                                             
                tmr_registers(1)(875)    <= not(global_tmr_voter(1)(874));                                                             
                tmr_registers(2)(875)    <= not(global_tmr_voter(2)(874));                                                             
 
                tmr_registers(0)(876)    <= not(global_tmr_voter(0)(875));                                                             
                tmr_registers(1)(876)    <= not(global_tmr_voter(1)(875));                                                             
                tmr_registers(2)(876)    <= not(global_tmr_voter(2)(875));                                                             
 
                tmr_registers(0)(877)    <= not(global_tmr_voter(0)(876));                                                             
                tmr_registers(1)(877)    <= not(global_tmr_voter(1)(876));                                                             
                tmr_registers(2)(877)    <= not(global_tmr_voter(2)(876));                                                             
 
                tmr_registers(0)(878)    <= not(global_tmr_voter(0)(877));                                                             
                tmr_registers(1)(878)    <= not(global_tmr_voter(1)(877));                                                             
                tmr_registers(2)(878)    <= not(global_tmr_voter(2)(877));                                                             
 
                tmr_registers(0)(879)    <= not(global_tmr_voter(0)(878));                                                             
                tmr_registers(1)(879)    <= not(global_tmr_voter(1)(878));                                                             
                tmr_registers(2)(879)    <= not(global_tmr_voter(2)(878));                                                             
 
                tmr_registers(0)(880)    <= not(global_tmr_voter(0)(879));                                                             
                tmr_registers(1)(880)    <= not(global_tmr_voter(1)(879));                                                             
                tmr_registers(2)(880)    <= not(global_tmr_voter(2)(879));                                                             
 
                tmr_registers(0)(881)    <= not(global_tmr_voter(0)(880));                                                             
                tmr_registers(1)(881)    <= not(global_tmr_voter(1)(880));                                                             
                tmr_registers(2)(881)    <= not(global_tmr_voter(2)(880));                                                             
 
                tmr_registers(0)(882)    <= not(global_tmr_voter(0)(881));                                                             
                tmr_registers(1)(882)    <= not(global_tmr_voter(1)(881));                                                             
                tmr_registers(2)(882)    <= not(global_tmr_voter(2)(881));                                                             
 
                tmr_registers(0)(883)    <= not(global_tmr_voter(0)(882));                                                             
                tmr_registers(1)(883)    <= not(global_tmr_voter(1)(882));                                                             
                tmr_registers(2)(883)    <= not(global_tmr_voter(2)(882));                                                             
 
                tmr_registers(0)(884)    <= not(global_tmr_voter(0)(883));                                                             
                tmr_registers(1)(884)    <= not(global_tmr_voter(1)(883));                                                             
                tmr_registers(2)(884)    <= not(global_tmr_voter(2)(883));                                                             
 
                tmr_registers(0)(885)    <= not(global_tmr_voter(0)(884));                                                             
                tmr_registers(1)(885)    <= not(global_tmr_voter(1)(884));                                                             
                tmr_registers(2)(885)    <= not(global_tmr_voter(2)(884));                                                             
 
                tmr_registers(0)(886)    <= not(global_tmr_voter(0)(885));                                                             
                tmr_registers(1)(886)    <= not(global_tmr_voter(1)(885));                                                             
                tmr_registers(2)(886)    <= not(global_tmr_voter(2)(885));                                                             
 
                tmr_registers(0)(887)    <= not(global_tmr_voter(0)(886));                                                             
                tmr_registers(1)(887)    <= not(global_tmr_voter(1)(886));                                                             
                tmr_registers(2)(887)    <= not(global_tmr_voter(2)(886));                                                             
 
                tmr_registers(0)(888)    <= not(global_tmr_voter(0)(887));                                                             
                tmr_registers(1)(888)    <= not(global_tmr_voter(1)(887));                                                             
                tmr_registers(2)(888)    <= not(global_tmr_voter(2)(887));                                                             
 
                tmr_registers(0)(889)    <= not(global_tmr_voter(0)(888));                                                             
                tmr_registers(1)(889)    <= not(global_tmr_voter(1)(888));                                                             
                tmr_registers(2)(889)    <= not(global_tmr_voter(2)(888));                                                             
 
                tmr_registers(0)(890)    <= not(global_tmr_voter(0)(889));                                                             
                tmr_registers(1)(890)    <= not(global_tmr_voter(1)(889));                                                             
                tmr_registers(2)(890)    <= not(global_tmr_voter(2)(889));                                                             
 
                tmr_registers(0)(891)    <= not(global_tmr_voter(0)(890));                                                             
                tmr_registers(1)(891)    <= not(global_tmr_voter(1)(890));                                                             
                tmr_registers(2)(891)    <= not(global_tmr_voter(2)(890));                                                             
 
                tmr_registers(0)(892)    <= not(global_tmr_voter(0)(891));                                                             
                tmr_registers(1)(892)    <= not(global_tmr_voter(1)(891));                                                             
                tmr_registers(2)(892)    <= not(global_tmr_voter(2)(891));                                                             
 
                tmr_registers(0)(893)    <= not(global_tmr_voter(0)(892));                                                             
                tmr_registers(1)(893)    <= not(global_tmr_voter(1)(892));                                                             
                tmr_registers(2)(893)    <= not(global_tmr_voter(2)(892));                                                             
 
                tmr_registers(0)(894)    <= not(global_tmr_voter(0)(893));                                                             
                tmr_registers(1)(894)    <= not(global_tmr_voter(1)(893));                                                             
                tmr_registers(2)(894)    <= not(global_tmr_voter(2)(893));                                                             
 
                tmr_registers(0)(895)    <= not(global_tmr_voter(0)(894));                                                             
                tmr_registers(1)(895)    <= not(global_tmr_voter(1)(894));                                                             
                tmr_registers(2)(895)    <= not(global_tmr_voter(2)(894));                                                             
 
                tmr_registers(0)(896)    <= not(global_tmr_voter(0)(895));                                                             
                tmr_registers(1)(896)    <= not(global_tmr_voter(1)(895));                                                             
                tmr_registers(2)(896)    <= not(global_tmr_voter(2)(895));                                                             
 
                tmr_registers(0)(897)    <= not(global_tmr_voter(0)(896));                                                             
                tmr_registers(1)(897)    <= not(global_tmr_voter(1)(896));                                                             
                tmr_registers(2)(897)    <= not(global_tmr_voter(2)(896));                                                             
 
                tmr_registers(0)(898)    <= not(global_tmr_voter(0)(897));                                                             
                tmr_registers(1)(898)    <= not(global_tmr_voter(1)(897));                                                             
                tmr_registers(2)(898)    <= not(global_tmr_voter(2)(897));                                                             
 
                tmr_registers(0)(899)    <= not(global_tmr_voter(0)(898));                                                             
                tmr_registers(1)(899)    <= not(global_tmr_voter(1)(898));                                                             
                tmr_registers(2)(899)    <= not(global_tmr_voter(2)(898));                                                             
 
                tmr_registers(0)(900)    <= not(global_tmr_voter(0)(899));                                                             
                tmr_registers(1)(900)    <= not(global_tmr_voter(1)(899));                                                             
                tmr_registers(2)(900)    <= not(global_tmr_voter(2)(899));                                                             
 
                tmr_registers(0)(901)    <= not(global_tmr_voter(0)(900));                                                             
                tmr_registers(1)(901)    <= not(global_tmr_voter(1)(900));                                                             
                tmr_registers(2)(901)    <= not(global_tmr_voter(2)(900));                                                             
 
                tmr_registers(0)(902)    <= not(global_tmr_voter(0)(901));                                                             
                tmr_registers(1)(902)    <= not(global_tmr_voter(1)(901));                                                             
                tmr_registers(2)(902)    <= not(global_tmr_voter(2)(901));                                                             
 
                tmr_registers(0)(903)    <= not(global_tmr_voter(0)(902));                                                             
                tmr_registers(1)(903)    <= not(global_tmr_voter(1)(902));                                                             
                tmr_registers(2)(903)    <= not(global_tmr_voter(2)(902));                                                             
 
                tmr_registers(0)(904)    <= not(global_tmr_voter(0)(903));                                                             
                tmr_registers(1)(904)    <= not(global_tmr_voter(1)(903));                                                             
                tmr_registers(2)(904)    <= not(global_tmr_voter(2)(903));                                                             
 
                tmr_registers(0)(905)    <= not(global_tmr_voter(0)(904));                                                             
                tmr_registers(1)(905)    <= not(global_tmr_voter(1)(904));                                                             
                tmr_registers(2)(905)    <= not(global_tmr_voter(2)(904));                                                             
 
                tmr_registers(0)(906)    <= not(global_tmr_voter(0)(905));                                                             
                tmr_registers(1)(906)    <= not(global_tmr_voter(1)(905));                                                             
                tmr_registers(2)(906)    <= not(global_tmr_voter(2)(905));                                                             
 
                tmr_registers(0)(907)    <= not(global_tmr_voter(0)(906));                                                             
                tmr_registers(1)(907)    <= not(global_tmr_voter(1)(906));                                                             
                tmr_registers(2)(907)    <= not(global_tmr_voter(2)(906));                                                             
 
                tmr_registers(0)(908)    <= not(global_tmr_voter(0)(907));                                                             
                tmr_registers(1)(908)    <= not(global_tmr_voter(1)(907));                                                             
                tmr_registers(2)(908)    <= not(global_tmr_voter(2)(907));                                                             
 
                tmr_registers(0)(909)    <= not(global_tmr_voter(0)(908));                                                             
                tmr_registers(1)(909)    <= not(global_tmr_voter(1)(908));                                                             
                tmr_registers(2)(909)    <= not(global_tmr_voter(2)(908));                                                             
 
                tmr_registers(0)(910)    <= not(global_tmr_voter(0)(909));                                                             
                tmr_registers(1)(910)    <= not(global_tmr_voter(1)(909));                                                             
                tmr_registers(2)(910)    <= not(global_tmr_voter(2)(909));                                                             
 
                tmr_registers(0)(911)    <= not(global_tmr_voter(0)(910));                                                             
                tmr_registers(1)(911)    <= not(global_tmr_voter(1)(910));                                                             
                tmr_registers(2)(911)    <= not(global_tmr_voter(2)(910));                                                             
 
                tmr_registers(0)(912)    <= not(global_tmr_voter(0)(911));                                                             
                tmr_registers(1)(912)    <= not(global_tmr_voter(1)(911));                                                             
                tmr_registers(2)(912)    <= not(global_tmr_voter(2)(911));                                                             
 
                tmr_registers(0)(913)    <= not(global_tmr_voter(0)(912));                                                             
                tmr_registers(1)(913)    <= not(global_tmr_voter(1)(912));                                                             
                tmr_registers(2)(913)    <= not(global_tmr_voter(2)(912));                                                             
 
                tmr_registers(0)(914)    <= not(global_tmr_voter(0)(913));                                                             
                tmr_registers(1)(914)    <= not(global_tmr_voter(1)(913));                                                             
                tmr_registers(2)(914)    <= not(global_tmr_voter(2)(913));                                                             
 
                tmr_registers(0)(915)    <= not(global_tmr_voter(0)(914));                                                             
                tmr_registers(1)(915)    <= not(global_tmr_voter(1)(914));                                                             
                tmr_registers(2)(915)    <= not(global_tmr_voter(2)(914));                                                             
 
                tmr_registers(0)(916)    <= not(global_tmr_voter(0)(915));                                                             
                tmr_registers(1)(916)    <= not(global_tmr_voter(1)(915));                                                             
                tmr_registers(2)(916)    <= not(global_tmr_voter(2)(915));                                                             
 
                tmr_registers(0)(917)    <= not(global_tmr_voter(0)(916));                                                             
                tmr_registers(1)(917)    <= not(global_tmr_voter(1)(916));                                                             
                tmr_registers(2)(917)    <= not(global_tmr_voter(2)(916));                                                             
 
                tmr_registers(0)(918)    <= not(global_tmr_voter(0)(917));                                                             
                tmr_registers(1)(918)    <= not(global_tmr_voter(1)(917));                                                             
                tmr_registers(2)(918)    <= not(global_tmr_voter(2)(917));                                                             
 
                tmr_registers(0)(919)    <= not(global_tmr_voter(0)(918));                                                             
                tmr_registers(1)(919)    <= not(global_tmr_voter(1)(918));                                                             
                tmr_registers(2)(919)    <= not(global_tmr_voter(2)(918));                                                             
 
                tmr_registers(0)(920)    <= not(global_tmr_voter(0)(919));                                                             
                tmr_registers(1)(920)    <= not(global_tmr_voter(1)(919));                                                             
                tmr_registers(2)(920)    <= not(global_tmr_voter(2)(919));                                                             
 
                tmr_registers(0)(921)    <= not(global_tmr_voter(0)(920));                                                             
                tmr_registers(1)(921)    <= not(global_tmr_voter(1)(920));                                                             
                tmr_registers(2)(921)    <= not(global_tmr_voter(2)(920));                                                             
 
                tmr_registers(0)(922)    <= not(global_tmr_voter(0)(921));                                                             
                tmr_registers(1)(922)    <= not(global_tmr_voter(1)(921));                                                             
                tmr_registers(2)(922)    <= not(global_tmr_voter(2)(921));                                                             
 
                tmr_registers(0)(923)    <= not(global_tmr_voter(0)(922));                                                             
                tmr_registers(1)(923)    <= not(global_tmr_voter(1)(922));                                                             
                tmr_registers(2)(923)    <= not(global_tmr_voter(2)(922));                                                             
 
                tmr_registers(0)(924)    <= not(global_tmr_voter(0)(923));                                                             
                tmr_registers(1)(924)    <= not(global_tmr_voter(1)(923));                                                             
                tmr_registers(2)(924)    <= not(global_tmr_voter(2)(923));                                                             
 
                tmr_registers(0)(925)    <= not(global_tmr_voter(0)(924));                                                             
                tmr_registers(1)(925)    <= not(global_tmr_voter(1)(924));                                                             
                tmr_registers(2)(925)    <= not(global_tmr_voter(2)(924));                                                             
 
                tmr_registers(0)(926)    <= not(global_tmr_voter(0)(925));                                                             
                tmr_registers(1)(926)    <= not(global_tmr_voter(1)(925));                                                             
                tmr_registers(2)(926)    <= not(global_tmr_voter(2)(925));                                                             
 
                tmr_registers(0)(927)    <= not(global_tmr_voter(0)(926));                                                             
                tmr_registers(1)(927)    <= not(global_tmr_voter(1)(926));                                                             
                tmr_registers(2)(927)    <= not(global_tmr_voter(2)(926));                                                             
 
                tmr_registers(0)(928)    <= not(global_tmr_voter(0)(927));                                                             
                tmr_registers(1)(928)    <= not(global_tmr_voter(1)(927));                                                             
                tmr_registers(2)(928)    <= not(global_tmr_voter(2)(927));                                                             
 
                tmr_registers(0)(929)    <= not(global_tmr_voter(0)(928));                                                             
                tmr_registers(1)(929)    <= not(global_tmr_voter(1)(928));                                                             
                tmr_registers(2)(929)    <= not(global_tmr_voter(2)(928));                                                             
 
                tmr_registers(0)(930)    <= not(global_tmr_voter(0)(929));                                                             
                tmr_registers(1)(930)    <= not(global_tmr_voter(1)(929));                                                             
                tmr_registers(2)(930)    <= not(global_tmr_voter(2)(929));                                                             
 
                tmr_registers(0)(931)    <= not(global_tmr_voter(0)(930));                                                             
                tmr_registers(1)(931)    <= not(global_tmr_voter(1)(930));                                                             
                tmr_registers(2)(931)    <= not(global_tmr_voter(2)(930));                                                             
 
                tmr_registers(0)(932)    <= not(global_tmr_voter(0)(931));                                                             
                tmr_registers(1)(932)    <= not(global_tmr_voter(1)(931));                                                             
                tmr_registers(2)(932)    <= not(global_tmr_voter(2)(931));                                                             
 
                tmr_registers(0)(933)    <= not(global_tmr_voter(0)(932));                                                             
                tmr_registers(1)(933)    <= not(global_tmr_voter(1)(932));                                                             
                tmr_registers(2)(933)    <= not(global_tmr_voter(2)(932));                                                             
 
                tmr_registers(0)(934)    <= not(global_tmr_voter(0)(933));                                                             
                tmr_registers(1)(934)    <= not(global_tmr_voter(1)(933));                                                             
                tmr_registers(2)(934)    <= not(global_tmr_voter(2)(933));                                                             
 
                tmr_registers(0)(935)    <= not(global_tmr_voter(0)(934));                                                             
                tmr_registers(1)(935)    <= not(global_tmr_voter(1)(934));                                                             
                tmr_registers(2)(935)    <= not(global_tmr_voter(2)(934));                                                             
 
                tmr_registers(0)(936)    <= not(global_tmr_voter(0)(935));                                                             
                tmr_registers(1)(936)    <= not(global_tmr_voter(1)(935));                                                             
                tmr_registers(2)(936)    <= not(global_tmr_voter(2)(935));                                                             
 
                tmr_registers(0)(937)    <= not(global_tmr_voter(0)(936));                                                             
                tmr_registers(1)(937)    <= not(global_tmr_voter(1)(936));                                                             
                tmr_registers(2)(937)    <= not(global_tmr_voter(2)(936));                                                             
 
                tmr_registers(0)(938)    <= not(global_tmr_voter(0)(937));                                                             
                tmr_registers(1)(938)    <= not(global_tmr_voter(1)(937));                                                             
                tmr_registers(2)(938)    <= not(global_tmr_voter(2)(937));                                                             
 
                tmr_registers(0)(939)    <= not(global_tmr_voter(0)(938));                                                             
                tmr_registers(1)(939)    <= not(global_tmr_voter(1)(938));                                                             
                tmr_registers(2)(939)    <= not(global_tmr_voter(2)(938));                                                             
 
                tmr_registers(0)(940)    <= not(global_tmr_voter(0)(939));                                                             
                tmr_registers(1)(940)    <= not(global_tmr_voter(1)(939));                                                             
                tmr_registers(2)(940)    <= not(global_tmr_voter(2)(939));                                                             
 
                tmr_registers(0)(941)    <= not(global_tmr_voter(0)(940));                                                             
                tmr_registers(1)(941)    <= not(global_tmr_voter(1)(940));                                                             
                tmr_registers(2)(941)    <= not(global_tmr_voter(2)(940));                                                             
 
                tmr_registers(0)(942)    <= not(global_tmr_voter(0)(941));                                                             
                tmr_registers(1)(942)    <= not(global_tmr_voter(1)(941));                                                             
                tmr_registers(2)(942)    <= not(global_tmr_voter(2)(941));                                                             
 
                tmr_registers(0)(943)    <= not(global_tmr_voter(0)(942));                                                             
                tmr_registers(1)(943)    <= not(global_tmr_voter(1)(942));                                                             
                tmr_registers(2)(943)    <= not(global_tmr_voter(2)(942));                                                             
 
                tmr_registers(0)(944)    <= not(global_tmr_voter(0)(943));                                                             
                tmr_registers(1)(944)    <= not(global_tmr_voter(1)(943));                                                             
                tmr_registers(2)(944)    <= not(global_tmr_voter(2)(943));                                                             
 
                tmr_registers(0)(945)    <= not(global_tmr_voter(0)(944));                                                             
                tmr_registers(1)(945)    <= not(global_tmr_voter(1)(944));                                                             
                tmr_registers(2)(945)    <= not(global_tmr_voter(2)(944));                                                             
 
                tmr_registers(0)(946)    <= not(global_tmr_voter(0)(945));                                                             
                tmr_registers(1)(946)    <= not(global_tmr_voter(1)(945));                                                             
                tmr_registers(2)(946)    <= not(global_tmr_voter(2)(945));                                                             
 
                tmr_registers(0)(947)    <= not(global_tmr_voter(0)(946));                                                             
                tmr_registers(1)(947)    <= not(global_tmr_voter(1)(946));                                                             
                tmr_registers(2)(947)    <= not(global_tmr_voter(2)(946));                                                             
 
                tmr_registers(0)(948)    <= not(global_tmr_voter(0)(947));                                                             
                tmr_registers(1)(948)    <= not(global_tmr_voter(1)(947));                                                             
                tmr_registers(2)(948)    <= not(global_tmr_voter(2)(947));                                                             
 
                tmr_registers(0)(949)    <= not(global_tmr_voter(0)(948));                                                             
                tmr_registers(1)(949)    <= not(global_tmr_voter(1)(948));                                                             
                tmr_registers(2)(949)    <= not(global_tmr_voter(2)(948));                                                             
 
                tmr_registers(0)(950)    <= not(global_tmr_voter(0)(949));                                                             
                tmr_registers(1)(950)    <= not(global_tmr_voter(1)(949));                                                             
                tmr_registers(2)(950)    <= not(global_tmr_voter(2)(949));                                                             
 
                tmr_registers(0)(951)    <= not(global_tmr_voter(0)(950));                                                             
                tmr_registers(1)(951)    <= not(global_tmr_voter(1)(950));                                                             
                tmr_registers(2)(951)    <= not(global_tmr_voter(2)(950));                                                             
 
                tmr_registers(0)(952)    <= not(global_tmr_voter(0)(951));                                                             
                tmr_registers(1)(952)    <= not(global_tmr_voter(1)(951));                                                             
                tmr_registers(2)(952)    <= not(global_tmr_voter(2)(951));                                                             
 
                tmr_registers(0)(953)    <= not(global_tmr_voter(0)(952));                                                             
                tmr_registers(1)(953)    <= not(global_tmr_voter(1)(952));                                                             
                tmr_registers(2)(953)    <= not(global_tmr_voter(2)(952));                                                             
 
                tmr_registers(0)(954)    <= not(global_tmr_voter(0)(953));                                                             
                tmr_registers(1)(954)    <= not(global_tmr_voter(1)(953));                                                             
                tmr_registers(2)(954)    <= not(global_tmr_voter(2)(953));                                                             
 
                tmr_registers(0)(955)    <= not(global_tmr_voter(0)(954));                                                             
                tmr_registers(1)(955)    <= not(global_tmr_voter(1)(954));                                                             
                tmr_registers(2)(955)    <= not(global_tmr_voter(2)(954));                                                             
 
                tmr_registers(0)(956)    <= not(global_tmr_voter(0)(955));                                                             
                tmr_registers(1)(956)    <= not(global_tmr_voter(1)(955));                                                             
                tmr_registers(2)(956)    <= not(global_tmr_voter(2)(955));                                                             
 
                tmr_registers(0)(957)    <= not(global_tmr_voter(0)(956));                                                             
                tmr_registers(1)(957)    <= not(global_tmr_voter(1)(956));                                                             
                tmr_registers(2)(957)    <= not(global_tmr_voter(2)(956));                                                             
 
                tmr_registers(0)(958)    <= not(global_tmr_voter(0)(957));                                                             
                tmr_registers(1)(958)    <= not(global_tmr_voter(1)(957));                                                             
                tmr_registers(2)(958)    <= not(global_tmr_voter(2)(957));                                                             
 
                tmr_registers(0)(959)    <= not(global_tmr_voter(0)(958));                                                             
                tmr_registers(1)(959)    <= not(global_tmr_voter(1)(958));                                                             
                tmr_registers(2)(959)    <= not(global_tmr_voter(2)(958));                                                             
 
                tmr_registers(0)(960)    <= not(global_tmr_voter(0)(959));                                                             
                tmr_registers(1)(960)    <= not(global_tmr_voter(1)(959));                                                             
                tmr_registers(2)(960)    <= not(global_tmr_voter(2)(959));                                                             
 
                tmr_registers(0)(961)    <= not(global_tmr_voter(0)(960));                                                             
                tmr_registers(1)(961)    <= not(global_tmr_voter(1)(960));                                                             
                tmr_registers(2)(961)    <= not(global_tmr_voter(2)(960));                                                             
 
                tmr_registers(0)(962)    <= not(global_tmr_voter(0)(961));                                                             
                tmr_registers(1)(962)    <= not(global_tmr_voter(1)(961));                                                             
                tmr_registers(2)(962)    <= not(global_tmr_voter(2)(961));                                                             
 
                tmr_registers(0)(963)    <= not(global_tmr_voter(0)(962));                                                             
                tmr_registers(1)(963)    <= not(global_tmr_voter(1)(962));                                                             
                tmr_registers(2)(963)    <= not(global_tmr_voter(2)(962));                                                             
 
                tmr_registers(0)(964)    <= not(global_tmr_voter(0)(963));                                                             
                tmr_registers(1)(964)    <= not(global_tmr_voter(1)(963));                                                             
                tmr_registers(2)(964)    <= not(global_tmr_voter(2)(963));                                                             
 
                tmr_registers(0)(965)    <= not(global_tmr_voter(0)(964));                                                             
                tmr_registers(1)(965)    <= not(global_tmr_voter(1)(964));                                                             
                tmr_registers(2)(965)    <= not(global_tmr_voter(2)(964));                                                             
 
                tmr_registers(0)(966)    <= not(global_tmr_voter(0)(965));                                                             
                tmr_registers(1)(966)    <= not(global_tmr_voter(1)(965));                                                             
                tmr_registers(2)(966)    <= not(global_tmr_voter(2)(965));                                                             
 
                tmr_registers(0)(967)    <= not(global_tmr_voter(0)(966));                                                             
                tmr_registers(1)(967)    <= not(global_tmr_voter(1)(966));                                                             
                tmr_registers(2)(967)    <= not(global_tmr_voter(2)(966));                                                             
 
                tmr_registers(0)(968)    <= not(global_tmr_voter(0)(967));                                                             
                tmr_registers(1)(968)    <= not(global_tmr_voter(1)(967));                                                             
                tmr_registers(2)(968)    <= not(global_tmr_voter(2)(967));                                                             
 
                tmr_registers(0)(969)    <= not(global_tmr_voter(0)(968));                                                             
                tmr_registers(1)(969)    <= not(global_tmr_voter(1)(968));                                                             
                tmr_registers(2)(969)    <= not(global_tmr_voter(2)(968));                                                             
 
                tmr_registers(0)(970)    <= not(global_tmr_voter(0)(969));                                                             
                tmr_registers(1)(970)    <= not(global_tmr_voter(1)(969));                                                             
                tmr_registers(2)(970)    <= not(global_tmr_voter(2)(969));                                                             
 
                tmr_registers(0)(971)    <= not(global_tmr_voter(0)(970));                                                             
                tmr_registers(1)(971)    <= not(global_tmr_voter(1)(970));                                                             
                tmr_registers(2)(971)    <= not(global_tmr_voter(2)(970));                                                             
 
                tmr_registers(0)(972)    <= not(global_tmr_voter(0)(971));                                                             
                tmr_registers(1)(972)    <= not(global_tmr_voter(1)(971));                                                             
                tmr_registers(2)(972)    <= not(global_tmr_voter(2)(971));                                                             
 
                tmr_registers(0)(973)    <= not(global_tmr_voter(0)(972));                                                             
                tmr_registers(1)(973)    <= not(global_tmr_voter(1)(972));                                                             
                tmr_registers(2)(973)    <= not(global_tmr_voter(2)(972));                                                             
 
                tmr_registers(0)(974)    <= not(global_tmr_voter(0)(973));                                                             
                tmr_registers(1)(974)    <= not(global_tmr_voter(1)(973));                                                             
                tmr_registers(2)(974)    <= not(global_tmr_voter(2)(973));                                                             
 
                tmr_registers(0)(975)    <= not(global_tmr_voter(0)(974));                                                             
                tmr_registers(1)(975)    <= not(global_tmr_voter(1)(974));                                                             
                tmr_registers(2)(975)    <= not(global_tmr_voter(2)(974));                                                             
 
                tmr_registers(0)(976)    <= not(global_tmr_voter(0)(975));                                                             
                tmr_registers(1)(976)    <= not(global_tmr_voter(1)(975));                                                             
                tmr_registers(2)(976)    <= not(global_tmr_voter(2)(975));                                                             
 
                tmr_registers(0)(977)    <= not(global_tmr_voter(0)(976));                                                             
                tmr_registers(1)(977)    <= not(global_tmr_voter(1)(976));                                                             
                tmr_registers(2)(977)    <= not(global_tmr_voter(2)(976));                                                             
 
                tmr_registers(0)(978)    <= not(global_tmr_voter(0)(977));                                                             
                tmr_registers(1)(978)    <= not(global_tmr_voter(1)(977));                                                             
                tmr_registers(2)(978)    <= not(global_tmr_voter(2)(977));                                                             
 
                tmr_registers(0)(979)    <= not(global_tmr_voter(0)(978));                                                             
                tmr_registers(1)(979)    <= not(global_tmr_voter(1)(978));                                                             
                tmr_registers(2)(979)    <= not(global_tmr_voter(2)(978));                                                             
 
                tmr_registers(0)(980)    <= not(global_tmr_voter(0)(979));                                                             
                tmr_registers(1)(980)    <= not(global_tmr_voter(1)(979));                                                             
                tmr_registers(2)(980)    <= not(global_tmr_voter(2)(979));                                                             
 
                tmr_registers(0)(981)    <= not(global_tmr_voter(0)(980));                                                             
                tmr_registers(1)(981)    <= not(global_tmr_voter(1)(980));                                                             
                tmr_registers(2)(981)    <= not(global_tmr_voter(2)(980));                                                             
 
                tmr_registers(0)(982)    <= not(global_tmr_voter(0)(981));                                                             
                tmr_registers(1)(982)    <= not(global_tmr_voter(1)(981));                                                             
                tmr_registers(2)(982)    <= not(global_tmr_voter(2)(981));                                                             
 
                tmr_registers(0)(983)    <= not(global_tmr_voter(0)(982));                                                             
                tmr_registers(1)(983)    <= not(global_tmr_voter(1)(982));                                                             
                tmr_registers(2)(983)    <= not(global_tmr_voter(2)(982));                                                             
 
                tmr_registers(0)(984)    <= not(global_tmr_voter(0)(983));                                                             
                tmr_registers(1)(984)    <= not(global_tmr_voter(1)(983));                                                             
                tmr_registers(2)(984)    <= not(global_tmr_voter(2)(983));                                                             
 
                tmr_registers(0)(985)    <= not(global_tmr_voter(0)(984));                                                             
                tmr_registers(1)(985)    <= not(global_tmr_voter(1)(984));                                                             
                tmr_registers(2)(985)    <= not(global_tmr_voter(2)(984));                                                             
 
                tmr_registers(0)(986)    <= not(global_tmr_voter(0)(985));                                                             
                tmr_registers(1)(986)    <= not(global_tmr_voter(1)(985));                                                             
                tmr_registers(2)(986)    <= not(global_tmr_voter(2)(985));                                                             
 
                tmr_registers(0)(987)    <= not(global_tmr_voter(0)(986));                                                             
                tmr_registers(1)(987)    <= not(global_tmr_voter(1)(986));                                                             
                tmr_registers(2)(987)    <= not(global_tmr_voter(2)(986));                                                             
 
                tmr_registers(0)(988)    <= not(global_tmr_voter(0)(987));                                                             
                tmr_registers(1)(988)    <= not(global_tmr_voter(1)(987));                                                             
                tmr_registers(2)(988)    <= not(global_tmr_voter(2)(987));                                                             
 
                tmr_registers(0)(989)    <= not(global_tmr_voter(0)(988));                                                             
                tmr_registers(1)(989)    <= not(global_tmr_voter(1)(988));                                                             
                tmr_registers(2)(989)    <= not(global_tmr_voter(2)(988));                                                             
 
                tmr_registers(0)(990)    <= not(global_tmr_voter(0)(989));                                                             
                tmr_registers(1)(990)    <= not(global_tmr_voter(1)(989));                                                             
                tmr_registers(2)(990)    <= not(global_tmr_voter(2)(989));                                                             
 
                tmr_registers(0)(991)    <= not(global_tmr_voter(0)(990));                                                             
                tmr_registers(1)(991)    <= not(global_tmr_voter(1)(990));                                                             
                tmr_registers(2)(991)    <= not(global_tmr_voter(2)(990));                                                             
 
                tmr_registers(0)(992)    <= not(global_tmr_voter(0)(991));                                                             
                tmr_registers(1)(992)    <= not(global_tmr_voter(1)(991));                                                             
                tmr_registers(2)(992)    <= not(global_tmr_voter(2)(991));                                                             
 
                tmr_registers(0)(993)    <= not(global_tmr_voter(0)(992));                                                             
                tmr_registers(1)(993)    <= not(global_tmr_voter(1)(992));                                                             
                tmr_registers(2)(993)    <= not(global_tmr_voter(2)(992));                                                             
 
                tmr_registers(0)(994)    <= not(global_tmr_voter(0)(993));                                                             
                tmr_registers(1)(994)    <= not(global_tmr_voter(1)(993));                                                             
                tmr_registers(2)(994)    <= not(global_tmr_voter(2)(993));                                                             
 
                tmr_registers(0)(995)    <= not(global_tmr_voter(0)(994));                                                             
                tmr_registers(1)(995)    <= not(global_tmr_voter(1)(994));                                                             
                tmr_registers(2)(995)    <= not(global_tmr_voter(2)(994));                                                             
 
                tmr_registers(0)(996)    <= not(global_tmr_voter(0)(995));                                                             
                tmr_registers(1)(996)    <= not(global_tmr_voter(1)(995));                                                             
                tmr_registers(2)(996)    <= not(global_tmr_voter(2)(995));                                                             
 
                tmr_registers(0)(997)    <= not(global_tmr_voter(0)(996));                                                             
                tmr_registers(1)(997)    <= not(global_tmr_voter(1)(996));                                                             
                tmr_registers(2)(997)    <= not(global_tmr_voter(2)(996));                                                             
 
                tmr_registers(0)(998)    <= not(global_tmr_voter(0)(997));                                                             
                tmr_registers(1)(998)    <= not(global_tmr_voter(1)(997));                                                             
                tmr_registers(2)(998)    <= not(global_tmr_voter(2)(997));                                                             
 
                tmr_registers(0)(999)    <= not(global_tmr_voter(0)(998));                                                             
                tmr_registers(1)(999)    <= not(global_tmr_voter(1)(998));                                                             
                tmr_registers(2)(999)    <= not(global_tmr_voter(2)(998));                                                             
 
                                                                                                                                         
        end if;                                                                                                                          
    end process;                                                                                                                         
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Voter                                                                                                                             
    ------------------------------------------                                                                                           
                                                                                                                                         
        global_tmr_voter(0)(0)  <= data_in;                                                                                              
        global_tmr_voter(1)(0)  <= data_in;                                                                                              
        global_tmr_voter(2)(0)  <= data_in;                                                                                              
                                                                                                                                     
        global_tmr_voter(0)(1)  <=    (tmr_registers(0)(1) and tmr_registers(1)(1)) or                                            
                            (tmr_registers(1)(1) and tmr_registers(2)(1)) or                                                       
                            (tmr_registers(0)(1) and tmr_registers(2)(1));                                                         
                                                                                                                                     
        global_tmr_voter(0)(2)  <=    (tmr_registers(0)(2) and tmr_registers(1)(2)) or                                            
                            (tmr_registers(1)(2) and tmr_registers(2)(2)) or                                                       
                            (tmr_registers(0)(2) and tmr_registers(2)(2));                                                         
                                                                                                                                     
        global_tmr_voter(0)(3)  <=    (tmr_registers(0)(3) and tmr_registers(1)(3)) or                                            
                            (tmr_registers(1)(3) and tmr_registers(2)(3)) or                                                       
                            (tmr_registers(0)(3) and tmr_registers(2)(3));                                                         
                                                                                                                                     
        global_tmr_voter(0)(4)  <=    (tmr_registers(0)(4) and tmr_registers(1)(4)) or                                            
                            (tmr_registers(1)(4) and tmr_registers(2)(4)) or                                                       
                            (tmr_registers(0)(4) and tmr_registers(2)(4));                                                         
                                                                                                                                     
        global_tmr_voter(0)(5)  <=    (tmr_registers(0)(5) and tmr_registers(1)(5)) or                                            
                            (tmr_registers(1)(5) and tmr_registers(2)(5)) or                                                       
                            (tmr_registers(0)(5) and tmr_registers(2)(5));                                                         
                                                                                                                                     
        global_tmr_voter(0)(6)  <=    (tmr_registers(0)(6) and tmr_registers(1)(6)) or                                            
                            (tmr_registers(1)(6) and tmr_registers(2)(6)) or                                                       
                            (tmr_registers(0)(6) and tmr_registers(2)(6));                                                         
                                                                                                                                     
        global_tmr_voter(0)(7)  <=    (tmr_registers(0)(7) and tmr_registers(1)(7)) or                                            
                            (tmr_registers(1)(7) and tmr_registers(2)(7)) or                                                       
                            (tmr_registers(0)(7) and tmr_registers(2)(7));                                                         
                                                                                                                                     
        global_tmr_voter(0)(8)  <=    (tmr_registers(0)(8) and tmr_registers(1)(8)) or                                            
                            (tmr_registers(1)(8) and tmr_registers(2)(8)) or                                                       
                            (tmr_registers(0)(8) and tmr_registers(2)(8));                                                         
                                                                                                                                     
        global_tmr_voter(0)(9)  <=    (tmr_registers(0)(9) and tmr_registers(1)(9)) or                                            
                            (tmr_registers(1)(9) and tmr_registers(2)(9)) or                                                       
                            (tmr_registers(0)(9) and tmr_registers(2)(9));                                                         
                                                                                                                                     
        global_tmr_voter(0)(10)  <=    (tmr_registers(0)(10) and tmr_registers(1)(10)) or                                            
                            (tmr_registers(1)(10) and tmr_registers(2)(10)) or                                                       
                            (tmr_registers(0)(10) and tmr_registers(2)(10));                                                         
                                                                                                                                     
        global_tmr_voter(0)(11)  <=    (tmr_registers(0)(11) and tmr_registers(1)(11)) or                                            
                            (tmr_registers(1)(11) and tmr_registers(2)(11)) or                                                       
                            (tmr_registers(0)(11) and tmr_registers(2)(11));                                                         
                                                                                                                                     
        global_tmr_voter(0)(12)  <=    (tmr_registers(0)(12) and tmr_registers(1)(12)) or                                            
                            (tmr_registers(1)(12) and tmr_registers(2)(12)) or                                                       
                            (tmr_registers(0)(12) and tmr_registers(2)(12));                                                         
                                                                                                                                     
        global_tmr_voter(0)(13)  <=    (tmr_registers(0)(13) and tmr_registers(1)(13)) or                                            
                            (tmr_registers(1)(13) and tmr_registers(2)(13)) or                                                       
                            (tmr_registers(0)(13) and tmr_registers(2)(13));                                                         
                                                                                                                                     
        global_tmr_voter(0)(14)  <=    (tmr_registers(0)(14) and tmr_registers(1)(14)) or                                            
                            (tmr_registers(1)(14) and tmr_registers(2)(14)) or                                                       
                            (tmr_registers(0)(14) and tmr_registers(2)(14));                                                         
                                                                                                                                     
        global_tmr_voter(0)(15)  <=    (tmr_registers(0)(15) and tmr_registers(1)(15)) or                                            
                            (tmr_registers(1)(15) and tmr_registers(2)(15)) or                                                       
                            (tmr_registers(0)(15) and tmr_registers(2)(15));                                                         
                                                                                                                                     
        global_tmr_voter(0)(16)  <=    (tmr_registers(0)(16) and tmr_registers(1)(16)) or                                            
                            (tmr_registers(1)(16) and tmr_registers(2)(16)) or                                                       
                            (tmr_registers(0)(16) and tmr_registers(2)(16));                                                         
                                                                                                                                     
        global_tmr_voter(0)(17)  <=    (tmr_registers(0)(17) and tmr_registers(1)(17)) or                                            
                            (tmr_registers(1)(17) and tmr_registers(2)(17)) or                                                       
                            (tmr_registers(0)(17) and tmr_registers(2)(17));                                                         
                                                                                                                                     
        global_tmr_voter(0)(18)  <=    (tmr_registers(0)(18) and tmr_registers(1)(18)) or                                            
                            (tmr_registers(1)(18) and tmr_registers(2)(18)) or                                                       
                            (tmr_registers(0)(18) and tmr_registers(2)(18));                                                         
                                                                                                                                     
        global_tmr_voter(0)(19)  <=    (tmr_registers(0)(19) and tmr_registers(1)(19)) or                                            
                            (tmr_registers(1)(19) and tmr_registers(2)(19)) or                                                       
                            (tmr_registers(0)(19) and tmr_registers(2)(19));                                                         
                                                                                                                                     
        global_tmr_voter(0)(20)  <=    (tmr_registers(0)(20) and tmr_registers(1)(20)) or                                            
                            (tmr_registers(1)(20) and tmr_registers(2)(20)) or                                                       
                            (tmr_registers(0)(20) and tmr_registers(2)(20));                                                         
                                                                                                                                     
        global_tmr_voter(0)(21)  <=    (tmr_registers(0)(21) and tmr_registers(1)(21)) or                                            
                            (tmr_registers(1)(21) and tmr_registers(2)(21)) or                                                       
                            (tmr_registers(0)(21) and tmr_registers(2)(21));                                                         
                                                                                                                                     
        global_tmr_voter(0)(22)  <=    (tmr_registers(0)(22) and tmr_registers(1)(22)) or                                            
                            (tmr_registers(1)(22) and tmr_registers(2)(22)) or                                                       
                            (tmr_registers(0)(22) and tmr_registers(2)(22));                                                         
                                                                                                                                     
        global_tmr_voter(0)(23)  <=    (tmr_registers(0)(23) and tmr_registers(1)(23)) or                                            
                            (tmr_registers(1)(23) and tmr_registers(2)(23)) or                                                       
                            (tmr_registers(0)(23) and tmr_registers(2)(23));                                                         
                                                                                                                                     
        global_tmr_voter(0)(24)  <=    (tmr_registers(0)(24) and tmr_registers(1)(24)) or                                            
                            (tmr_registers(1)(24) and tmr_registers(2)(24)) or                                                       
                            (tmr_registers(0)(24) and tmr_registers(2)(24));                                                         
                                                                                                                                     
        global_tmr_voter(0)(25)  <=    (tmr_registers(0)(25) and tmr_registers(1)(25)) or                                            
                            (tmr_registers(1)(25) and tmr_registers(2)(25)) or                                                       
                            (tmr_registers(0)(25) and tmr_registers(2)(25));                                                         
                                                                                                                                     
        global_tmr_voter(0)(26)  <=    (tmr_registers(0)(26) and tmr_registers(1)(26)) or                                            
                            (tmr_registers(1)(26) and tmr_registers(2)(26)) or                                                       
                            (tmr_registers(0)(26) and tmr_registers(2)(26));                                                         
                                                                                                                                     
        global_tmr_voter(0)(27)  <=    (tmr_registers(0)(27) and tmr_registers(1)(27)) or                                            
                            (tmr_registers(1)(27) and tmr_registers(2)(27)) or                                                       
                            (tmr_registers(0)(27) and tmr_registers(2)(27));                                                         
                                                                                                                                     
        global_tmr_voter(0)(28)  <=    (tmr_registers(0)(28) and tmr_registers(1)(28)) or                                            
                            (tmr_registers(1)(28) and tmr_registers(2)(28)) or                                                       
                            (tmr_registers(0)(28) and tmr_registers(2)(28));                                                         
                                                                                                                                     
        global_tmr_voter(0)(29)  <=    (tmr_registers(0)(29) and tmr_registers(1)(29)) or                                            
                            (tmr_registers(1)(29) and tmr_registers(2)(29)) or                                                       
                            (tmr_registers(0)(29) and tmr_registers(2)(29));                                                         
                                                                                                                                     
        global_tmr_voter(0)(30)  <=    (tmr_registers(0)(30) and tmr_registers(1)(30)) or                                            
                            (tmr_registers(1)(30) and tmr_registers(2)(30)) or                                                       
                            (tmr_registers(0)(30) and tmr_registers(2)(30));                                                         
                                                                                                                                     
        global_tmr_voter(0)(31)  <=    (tmr_registers(0)(31) and tmr_registers(1)(31)) or                                            
                            (tmr_registers(1)(31) and tmr_registers(2)(31)) or                                                       
                            (tmr_registers(0)(31) and tmr_registers(2)(31));                                                         
                                                                                                                                     
        global_tmr_voter(0)(32)  <=    (tmr_registers(0)(32) and tmr_registers(1)(32)) or                                            
                            (tmr_registers(1)(32) and tmr_registers(2)(32)) or                                                       
                            (tmr_registers(0)(32) and tmr_registers(2)(32));                                                         
                                                                                                                                     
        global_tmr_voter(0)(33)  <=    (tmr_registers(0)(33) and tmr_registers(1)(33)) or                                            
                            (tmr_registers(1)(33) and tmr_registers(2)(33)) or                                                       
                            (tmr_registers(0)(33) and tmr_registers(2)(33));                                                         
                                                                                                                                     
        global_tmr_voter(0)(34)  <=    (tmr_registers(0)(34) and tmr_registers(1)(34)) or                                            
                            (tmr_registers(1)(34) and tmr_registers(2)(34)) or                                                       
                            (tmr_registers(0)(34) and tmr_registers(2)(34));                                                         
                                                                                                                                     
        global_tmr_voter(0)(35)  <=    (tmr_registers(0)(35) and tmr_registers(1)(35)) or                                            
                            (tmr_registers(1)(35) and tmr_registers(2)(35)) or                                                       
                            (tmr_registers(0)(35) and tmr_registers(2)(35));                                                         
                                                                                                                                     
        global_tmr_voter(0)(36)  <=    (tmr_registers(0)(36) and tmr_registers(1)(36)) or                                            
                            (tmr_registers(1)(36) and tmr_registers(2)(36)) or                                                       
                            (tmr_registers(0)(36) and tmr_registers(2)(36));                                                         
                                                                                                                                     
        global_tmr_voter(0)(37)  <=    (tmr_registers(0)(37) and tmr_registers(1)(37)) or                                            
                            (tmr_registers(1)(37) and tmr_registers(2)(37)) or                                                       
                            (tmr_registers(0)(37) and tmr_registers(2)(37));                                                         
                                                                                                                                     
        global_tmr_voter(0)(38)  <=    (tmr_registers(0)(38) and tmr_registers(1)(38)) or                                            
                            (tmr_registers(1)(38) and tmr_registers(2)(38)) or                                                       
                            (tmr_registers(0)(38) and tmr_registers(2)(38));                                                         
                                                                                                                                     
        global_tmr_voter(0)(39)  <=    (tmr_registers(0)(39) and tmr_registers(1)(39)) or                                            
                            (tmr_registers(1)(39) and tmr_registers(2)(39)) or                                                       
                            (tmr_registers(0)(39) and tmr_registers(2)(39));                                                         
                                                                                                                                     
        global_tmr_voter(0)(40)  <=    (tmr_registers(0)(40) and tmr_registers(1)(40)) or                                            
                            (tmr_registers(1)(40) and tmr_registers(2)(40)) or                                                       
                            (tmr_registers(0)(40) and tmr_registers(2)(40));                                                         
                                                                                                                                     
        global_tmr_voter(0)(41)  <=    (tmr_registers(0)(41) and tmr_registers(1)(41)) or                                            
                            (tmr_registers(1)(41) and tmr_registers(2)(41)) or                                                       
                            (tmr_registers(0)(41) and tmr_registers(2)(41));                                                         
                                                                                                                                     
        global_tmr_voter(0)(42)  <=    (tmr_registers(0)(42) and tmr_registers(1)(42)) or                                            
                            (tmr_registers(1)(42) and tmr_registers(2)(42)) or                                                       
                            (tmr_registers(0)(42) and tmr_registers(2)(42));                                                         
                                                                                                                                     
        global_tmr_voter(0)(43)  <=    (tmr_registers(0)(43) and tmr_registers(1)(43)) or                                            
                            (tmr_registers(1)(43) and tmr_registers(2)(43)) or                                                       
                            (tmr_registers(0)(43) and tmr_registers(2)(43));                                                         
                                                                                                                                     
        global_tmr_voter(0)(44)  <=    (tmr_registers(0)(44) and tmr_registers(1)(44)) or                                            
                            (tmr_registers(1)(44) and tmr_registers(2)(44)) or                                                       
                            (tmr_registers(0)(44) and tmr_registers(2)(44));                                                         
                                                                                                                                     
        global_tmr_voter(0)(45)  <=    (tmr_registers(0)(45) and tmr_registers(1)(45)) or                                            
                            (tmr_registers(1)(45) and tmr_registers(2)(45)) or                                                       
                            (tmr_registers(0)(45) and tmr_registers(2)(45));                                                         
                                                                                                                                     
        global_tmr_voter(0)(46)  <=    (tmr_registers(0)(46) and tmr_registers(1)(46)) or                                            
                            (tmr_registers(1)(46) and tmr_registers(2)(46)) or                                                       
                            (tmr_registers(0)(46) and tmr_registers(2)(46));                                                         
                                                                                                                                     
        global_tmr_voter(0)(47)  <=    (tmr_registers(0)(47) and tmr_registers(1)(47)) or                                            
                            (tmr_registers(1)(47) and tmr_registers(2)(47)) or                                                       
                            (tmr_registers(0)(47) and tmr_registers(2)(47));                                                         
                                                                                                                                     
        global_tmr_voter(0)(48)  <=    (tmr_registers(0)(48) and tmr_registers(1)(48)) or                                            
                            (tmr_registers(1)(48) and tmr_registers(2)(48)) or                                                       
                            (tmr_registers(0)(48) and tmr_registers(2)(48));                                                         
                                                                                                                                     
        global_tmr_voter(0)(49)  <=    (tmr_registers(0)(49) and tmr_registers(1)(49)) or                                            
                            (tmr_registers(1)(49) and tmr_registers(2)(49)) or                                                       
                            (tmr_registers(0)(49) and tmr_registers(2)(49));                                                         
                                                                                                                                     
        global_tmr_voter(0)(50)  <=    (tmr_registers(0)(50) and tmr_registers(1)(50)) or                                            
                            (tmr_registers(1)(50) and tmr_registers(2)(50)) or                                                       
                            (tmr_registers(0)(50) and tmr_registers(2)(50));                                                         
                                                                                                                                     
        global_tmr_voter(0)(51)  <=    (tmr_registers(0)(51) and tmr_registers(1)(51)) or                                            
                            (tmr_registers(1)(51) and tmr_registers(2)(51)) or                                                       
                            (tmr_registers(0)(51) and tmr_registers(2)(51));                                                         
                                                                                                                                     
        global_tmr_voter(0)(52)  <=    (tmr_registers(0)(52) and tmr_registers(1)(52)) or                                            
                            (tmr_registers(1)(52) and tmr_registers(2)(52)) or                                                       
                            (tmr_registers(0)(52) and tmr_registers(2)(52));                                                         
                                                                                                                                     
        global_tmr_voter(0)(53)  <=    (tmr_registers(0)(53) and tmr_registers(1)(53)) or                                            
                            (tmr_registers(1)(53) and tmr_registers(2)(53)) or                                                       
                            (tmr_registers(0)(53) and tmr_registers(2)(53));                                                         
                                                                                                                                     
        global_tmr_voter(0)(54)  <=    (tmr_registers(0)(54) and tmr_registers(1)(54)) or                                            
                            (tmr_registers(1)(54) and tmr_registers(2)(54)) or                                                       
                            (tmr_registers(0)(54) and tmr_registers(2)(54));                                                         
                                                                                                                                     
        global_tmr_voter(0)(55)  <=    (tmr_registers(0)(55) and tmr_registers(1)(55)) or                                            
                            (tmr_registers(1)(55) and tmr_registers(2)(55)) or                                                       
                            (tmr_registers(0)(55) and tmr_registers(2)(55));                                                         
                                                                                                                                     
        global_tmr_voter(0)(56)  <=    (tmr_registers(0)(56) and tmr_registers(1)(56)) or                                            
                            (tmr_registers(1)(56) and tmr_registers(2)(56)) or                                                       
                            (tmr_registers(0)(56) and tmr_registers(2)(56));                                                         
                                                                                                                                     
        global_tmr_voter(0)(57)  <=    (tmr_registers(0)(57) and tmr_registers(1)(57)) or                                            
                            (tmr_registers(1)(57) and tmr_registers(2)(57)) or                                                       
                            (tmr_registers(0)(57) and tmr_registers(2)(57));                                                         
                                                                                                                                     
        global_tmr_voter(0)(58)  <=    (tmr_registers(0)(58) and tmr_registers(1)(58)) or                                            
                            (tmr_registers(1)(58) and tmr_registers(2)(58)) or                                                       
                            (tmr_registers(0)(58) and tmr_registers(2)(58));                                                         
                                                                                                                                     
        global_tmr_voter(0)(59)  <=    (tmr_registers(0)(59) and tmr_registers(1)(59)) or                                            
                            (tmr_registers(1)(59) and tmr_registers(2)(59)) or                                                       
                            (tmr_registers(0)(59) and tmr_registers(2)(59));                                                         
                                                                                                                                     
        global_tmr_voter(0)(60)  <=    (tmr_registers(0)(60) and tmr_registers(1)(60)) or                                            
                            (tmr_registers(1)(60) and tmr_registers(2)(60)) or                                                       
                            (tmr_registers(0)(60) and tmr_registers(2)(60));                                                         
                                                                                                                                     
        global_tmr_voter(0)(61)  <=    (tmr_registers(0)(61) and tmr_registers(1)(61)) or                                            
                            (tmr_registers(1)(61) and tmr_registers(2)(61)) or                                                       
                            (tmr_registers(0)(61) and tmr_registers(2)(61));                                                         
                                                                                                                                     
        global_tmr_voter(0)(62)  <=    (tmr_registers(0)(62) and tmr_registers(1)(62)) or                                            
                            (tmr_registers(1)(62) and tmr_registers(2)(62)) or                                                       
                            (tmr_registers(0)(62) and tmr_registers(2)(62));                                                         
                                                                                                                                     
        global_tmr_voter(0)(63)  <=    (tmr_registers(0)(63) and tmr_registers(1)(63)) or                                            
                            (tmr_registers(1)(63) and tmr_registers(2)(63)) or                                                       
                            (tmr_registers(0)(63) and tmr_registers(2)(63));                                                         
                                                                                                                                     
        global_tmr_voter(0)(64)  <=    (tmr_registers(0)(64) and tmr_registers(1)(64)) or                                            
                            (tmr_registers(1)(64) and tmr_registers(2)(64)) or                                                       
                            (tmr_registers(0)(64) and tmr_registers(2)(64));                                                         
                                                                                                                                     
        global_tmr_voter(0)(65)  <=    (tmr_registers(0)(65) and tmr_registers(1)(65)) or                                            
                            (tmr_registers(1)(65) and tmr_registers(2)(65)) or                                                       
                            (tmr_registers(0)(65) and tmr_registers(2)(65));                                                         
                                                                                                                                     
        global_tmr_voter(0)(66)  <=    (tmr_registers(0)(66) and tmr_registers(1)(66)) or                                            
                            (tmr_registers(1)(66) and tmr_registers(2)(66)) or                                                       
                            (tmr_registers(0)(66) and tmr_registers(2)(66));                                                         
                                                                                                                                     
        global_tmr_voter(0)(67)  <=    (tmr_registers(0)(67) and tmr_registers(1)(67)) or                                            
                            (tmr_registers(1)(67) and tmr_registers(2)(67)) or                                                       
                            (tmr_registers(0)(67) and tmr_registers(2)(67));                                                         
                                                                                                                                     
        global_tmr_voter(0)(68)  <=    (tmr_registers(0)(68) and tmr_registers(1)(68)) or                                            
                            (tmr_registers(1)(68) and tmr_registers(2)(68)) or                                                       
                            (tmr_registers(0)(68) and tmr_registers(2)(68));                                                         
                                                                                                                                     
        global_tmr_voter(0)(69)  <=    (tmr_registers(0)(69) and tmr_registers(1)(69)) or                                            
                            (tmr_registers(1)(69) and tmr_registers(2)(69)) or                                                       
                            (tmr_registers(0)(69) and tmr_registers(2)(69));                                                         
                                                                                                                                     
        global_tmr_voter(0)(70)  <=    (tmr_registers(0)(70) and tmr_registers(1)(70)) or                                            
                            (tmr_registers(1)(70) and tmr_registers(2)(70)) or                                                       
                            (tmr_registers(0)(70) and tmr_registers(2)(70));                                                         
                                                                                                                                     
        global_tmr_voter(0)(71)  <=    (tmr_registers(0)(71) and tmr_registers(1)(71)) or                                            
                            (tmr_registers(1)(71) and tmr_registers(2)(71)) or                                                       
                            (tmr_registers(0)(71) and tmr_registers(2)(71));                                                         
                                                                                                                                     
        global_tmr_voter(0)(72)  <=    (tmr_registers(0)(72) and tmr_registers(1)(72)) or                                            
                            (tmr_registers(1)(72) and tmr_registers(2)(72)) or                                                       
                            (tmr_registers(0)(72) and tmr_registers(2)(72));                                                         
                                                                                                                                     
        global_tmr_voter(0)(73)  <=    (tmr_registers(0)(73) and tmr_registers(1)(73)) or                                            
                            (tmr_registers(1)(73) and tmr_registers(2)(73)) or                                                       
                            (tmr_registers(0)(73) and tmr_registers(2)(73));                                                         
                                                                                                                                     
        global_tmr_voter(0)(74)  <=    (tmr_registers(0)(74) and tmr_registers(1)(74)) or                                            
                            (tmr_registers(1)(74) and tmr_registers(2)(74)) or                                                       
                            (tmr_registers(0)(74) and tmr_registers(2)(74));                                                         
                                                                                                                                     
        global_tmr_voter(0)(75)  <=    (tmr_registers(0)(75) and tmr_registers(1)(75)) or                                            
                            (tmr_registers(1)(75) and tmr_registers(2)(75)) or                                                       
                            (tmr_registers(0)(75) and tmr_registers(2)(75));                                                         
                                                                                                                                     
        global_tmr_voter(0)(76)  <=    (tmr_registers(0)(76) and tmr_registers(1)(76)) or                                            
                            (tmr_registers(1)(76) and tmr_registers(2)(76)) or                                                       
                            (tmr_registers(0)(76) and tmr_registers(2)(76));                                                         
                                                                                                                                     
        global_tmr_voter(0)(77)  <=    (tmr_registers(0)(77) and tmr_registers(1)(77)) or                                            
                            (tmr_registers(1)(77) and tmr_registers(2)(77)) or                                                       
                            (tmr_registers(0)(77) and tmr_registers(2)(77));                                                         
                                                                                                                                     
        global_tmr_voter(0)(78)  <=    (tmr_registers(0)(78) and tmr_registers(1)(78)) or                                            
                            (tmr_registers(1)(78) and tmr_registers(2)(78)) or                                                       
                            (tmr_registers(0)(78) and tmr_registers(2)(78));                                                         
                                                                                                                                     
        global_tmr_voter(0)(79)  <=    (tmr_registers(0)(79) and tmr_registers(1)(79)) or                                            
                            (tmr_registers(1)(79) and tmr_registers(2)(79)) or                                                       
                            (tmr_registers(0)(79) and tmr_registers(2)(79));                                                         
                                                                                                                                     
        global_tmr_voter(0)(80)  <=    (tmr_registers(0)(80) and tmr_registers(1)(80)) or                                            
                            (tmr_registers(1)(80) and tmr_registers(2)(80)) or                                                       
                            (tmr_registers(0)(80) and tmr_registers(2)(80));                                                         
                                                                                                                                     
        global_tmr_voter(0)(81)  <=    (tmr_registers(0)(81) and tmr_registers(1)(81)) or                                            
                            (tmr_registers(1)(81) and tmr_registers(2)(81)) or                                                       
                            (tmr_registers(0)(81) and tmr_registers(2)(81));                                                         
                                                                                                                                     
        global_tmr_voter(0)(82)  <=    (tmr_registers(0)(82) and tmr_registers(1)(82)) or                                            
                            (tmr_registers(1)(82) and tmr_registers(2)(82)) or                                                       
                            (tmr_registers(0)(82) and tmr_registers(2)(82));                                                         
                                                                                                                                     
        global_tmr_voter(0)(83)  <=    (tmr_registers(0)(83) and tmr_registers(1)(83)) or                                            
                            (tmr_registers(1)(83) and tmr_registers(2)(83)) or                                                       
                            (tmr_registers(0)(83) and tmr_registers(2)(83));                                                         
                                                                                                                                     
        global_tmr_voter(0)(84)  <=    (tmr_registers(0)(84) and tmr_registers(1)(84)) or                                            
                            (tmr_registers(1)(84) and tmr_registers(2)(84)) or                                                       
                            (tmr_registers(0)(84) and tmr_registers(2)(84));                                                         
                                                                                                                                     
        global_tmr_voter(0)(85)  <=    (tmr_registers(0)(85) and tmr_registers(1)(85)) or                                            
                            (tmr_registers(1)(85) and tmr_registers(2)(85)) or                                                       
                            (tmr_registers(0)(85) and tmr_registers(2)(85));                                                         
                                                                                                                                     
        global_tmr_voter(0)(86)  <=    (tmr_registers(0)(86) and tmr_registers(1)(86)) or                                            
                            (tmr_registers(1)(86) and tmr_registers(2)(86)) or                                                       
                            (tmr_registers(0)(86) and tmr_registers(2)(86));                                                         
                                                                                                                                     
        global_tmr_voter(0)(87)  <=    (tmr_registers(0)(87) and tmr_registers(1)(87)) or                                            
                            (tmr_registers(1)(87) and tmr_registers(2)(87)) or                                                       
                            (tmr_registers(0)(87) and tmr_registers(2)(87));                                                         
                                                                                                                                     
        global_tmr_voter(0)(88)  <=    (tmr_registers(0)(88) and tmr_registers(1)(88)) or                                            
                            (tmr_registers(1)(88) and tmr_registers(2)(88)) or                                                       
                            (tmr_registers(0)(88) and tmr_registers(2)(88));                                                         
                                                                                                                                     
        global_tmr_voter(0)(89)  <=    (tmr_registers(0)(89) and tmr_registers(1)(89)) or                                            
                            (tmr_registers(1)(89) and tmr_registers(2)(89)) or                                                       
                            (tmr_registers(0)(89) and tmr_registers(2)(89));                                                         
                                                                                                                                     
        global_tmr_voter(0)(90)  <=    (tmr_registers(0)(90) and tmr_registers(1)(90)) or                                            
                            (tmr_registers(1)(90) and tmr_registers(2)(90)) or                                                       
                            (tmr_registers(0)(90) and tmr_registers(2)(90));                                                         
                                                                                                                                     
        global_tmr_voter(0)(91)  <=    (tmr_registers(0)(91) and tmr_registers(1)(91)) or                                            
                            (tmr_registers(1)(91) and tmr_registers(2)(91)) or                                                       
                            (tmr_registers(0)(91) and tmr_registers(2)(91));                                                         
                                                                                                                                     
        global_tmr_voter(0)(92)  <=    (tmr_registers(0)(92) and tmr_registers(1)(92)) or                                            
                            (tmr_registers(1)(92) and tmr_registers(2)(92)) or                                                       
                            (tmr_registers(0)(92) and tmr_registers(2)(92));                                                         
                                                                                                                                     
        global_tmr_voter(0)(93)  <=    (tmr_registers(0)(93) and tmr_registers(1)(93)) or                                            
                            (tmr_registers(1)(93) and tmr_registers(2)(93)) or                                                       
                            (tmr_registers(0)(93) and tmr_registers(2)(93));                                                         
                                                                                                                                     
        global_tmr_voter(0)(94)  <=    (tmr_registers(0)(94) and tmr_registers(1)(94)) or                                            
                            (tmr_registers(1)(94) and tmr_registers(2)(94)) or                                                       
                            (tmr_registers(0)(94) and tmr_registers(2)(94));                                                         
                                                                                                                                     
        global_tmr_voter(0)(95)  <=    (tmr_registers(0)(95) and tmr_registers(1)(95)) or                                            
                            (tmr_registers(1)(95) and tmr_registers(2)(95)) or                                                       
                            (tmr_registers(0)(95) and tmr_registers(2)(95));                                                         
                                                                                                                                     
        global_tmr_voter(0)(96)  <=    (tmr_registers(0)(96) and tmr_registers(1)(96)) or                                            
                            (tmr_registers(1)(96) and tmr_registers(2)(96)) or                                                       
                            (tmr_registers(0)(96) and tmr_registers(2)(96));                                                         
                                                                                                                                     
        global_tmr_voter(0)(97)  <=    (tmr_registers(0)(97) and tmr_registers(1)(97)) or                                            
                            (tmr_registers(1)(97) and tmr_registers(2)(97)) or                                                       
                            (tmr_registers(0)(97) and tmr_registers(2)(97));                                                         
                                                                                                                                     
        global_tmr_voter(0)(98)  <=    (tmr_registers(0)(98) and tmr_registers(1)(98)) or                                            
                            (tmr_registers(1)(98) and tmr_registers(2)(98)) or                                                       
                            (tmr_registers(0)(98) and tmr_registers(2)(98));                                                         
                                                                                                                                     
        global_tmr_voter(0)(99)  <=    (tmr_registers(0)(99) and tmr_registers(1)(99)) or                                            
                            (tmr_registers(1)(99) and tmr_registers(2)(99)) or                                                       
                            (tmr_registers(0)(99) and tmr_registers(2)(99));                                                         
                                                                                                                                     
        global_tmr_voter(0)(100)  <=    (tmr_registers(0)(100) and tmr_registers(1)(100)) or                                            
                            (tmr_registers(1)(100) and tmr_registers(2)(100)) or                                                       
                            (tmr_registers(0)(100) and tmr_registers(2)(100));                                                         
                                                                                                                                     
        global_tmr_voter(0)(101)  <=    (tmr_registers(0)(101) and tmr_registers(1)(101)) or                                            
                            (tmr_registers(1)(101) and tmr_registers(2)(101)) or                                                       
                            (tmr_registers(0)(101) and tmr_registers(2)(101));                                                         
                                                                                                                                     
        global_tmr_voter(0)(102)  <=    (tmr_registers(0)(102) and tmr_registers(1)(102)) or                                            
                            (tmr_registers(1)(102) and tmr_registers(2)(102)) or                                                       
                            (tmr_registers(0)(102) and tmr_registers(2)(102));                                                         
                                                                                                                                     
        global_tmr_voter(0)(103)  <=    (tmr_registers(0)(103) and tmr_registers(1)(103)) or                                            
                            (tmr_registers(1)(103) and tmr_registers(2)(103)) or                                                       
                            (tmr_registers(0)(103) and tmr_registers(2)(103));                                                         
                                                                                                                                     
        global_tmr_voter(0)(104)  <=    (tmr_registers(0)(104) and tmr_registers(1)(104)) or                                            
                            (tmr_registers(1)(104) and tmr_registers(2)(104)) or                                                       
                            (tmr_registers(0)(104) and tmr_registers(2)(104));                                                         
                                                                                                                                     
        global_tmr_voter(0)(105)  <=    (tmr_registers(0)(105) and tmr_registers(1)(105)) or                                            
                            (tmr_registers(1)(105) and tmr_registers(2)(105)) or                                                       
                            (tmr_registers(0)(105) and tmr_registers(2)(105));                                                         
                                                                                                                                     
        global_tmr_voter(0)(106)  <=    (tmr_registers(0)(106) and tmr_registers(1)(106)) or                                            
                            (tmr_registers(1)(106) and tmr_registers(2)(106)) or                                                       
                            (tmr_registers(0)(106) and tmr_registers(2)(106));                                                         
                                                                                                                                     
        global_tmr_voter(0)(107)  <=    (tmr_registers(0)(107) and tmr_registers(1)(107)) or                                            
                            (tmr_registers(1)(107) and tmr_registers(2)(107)) or                                                       
                            (tmr_registers(0)(107) and tmr_registers(2)(107));                                                         
                                                                                                                                     
        global_tmr_voter(0)(108)  <=    (tmr_registers(0)(108) and tmr_registers(1)(108)) or                                            
                            (tmr_registers(1)(108) and tmr_registers(2)(108)) or                                                       
                            (tmr_registers(0)(108) and tmr_registers(2)(108));                                                         
                                                                                                                                     
        global_tmr_voter(0)(109)  <=    (tmr_registers(0)(109) and tmr_registers(1)(109)) or                                            
                            (tmr_registers(1)(109) and tmr_registers(2)(109)) or                                                       
                            (tmr_registers(0)(109) and tmr_registers(2)(109));                                                         
                                                                                                                                     
        global_tmr_voter(0)(110)  <=    (tmr_registers(0)(110) and tmr_registers(1)(110)) or                                            
                            (tmr_registers(1)(110) and tmr_registers(2)(110)) or                                                       
                            (tmr_registers(0)(110) and tmr_registers(2)(110));                                                         
                                                                                                                                     
        global_tmr_voter(0)(111)  <=    (tmr_registers(0)(111) and tmr_registers(1)(111)) or                                            
                            (tmr_registers(1)(111) and tmr_registers(2)(111)) or                                                       
                            (tmr_registers(0)(111) and tmr_registers(2)(111));                                                         
                                                                                                                                     
        global_tmr_voter(0)(112)  <=    (tmr_registers(0)(112) and tmr_registers(1)(112)) or                                            
                            (tmr_registers(1)(112) and tmr_registers(2)(112)) or                                                       
                            (tmr_registers(0)(112) and tmr_registers(2)(112));                                                         
                                                                                                                                     
        global_tmr_voter(0)(113)  <=    (tmr_registers(0)(113) and tmr_registers(1)(113)) or                                            
                            (tmr_registers(1)(113) and tmr_registers(2)(113)) or                                                       
                            (tmr_registers(0)(113) and tmr_registers(2)(113));                                                         
                                                                                                                                     
        global_tmr_voter(0)(114)  <=    (tmr_registers(0)(114) and tmr_registers(1)(114)) or                                            
                            (tmr_registers(1)(114) and tmr_registers(2)(114)) or                                                       
                            (tmr_registers(0)(114) and tmr_registers(2)(114));                                                         
                                                                                                                                     
        global_tmr_voter(0)(115)  <=    (tmr_registers(0)(115) and tmr_registers(1)(115)) or                                            
                            (tmr_registers(1)(115) and tmr_registers(2)(115)) or                                                       
                            (tmr_registers(0)(115) and tmr_registers(2)(115));                                                         
                                                                                                                                     
        global_tmr_voter(0)(116)  <=    (tmr_registers(0)(116) and tmr_registers(1)(116)) or                                            
                            (tmr_registers(1)(116) and tmr_registers(2)(116)) or                                                       
                            (tmr_registers(0)(116) and tmr_registers(2)(116));                                                         
                                                                                                                                     
        global_tmr_voter(0)(117)  <=    (tmr_registers(0)(117) and tmr_registers(1)(117)) or                                            
                            (tmr_registers(1)(117) and tmr_registers(2)(117)) or                                                       
                            (tmr_registers(0)(117) and tmr_registers(2)(117));                                                         
                                                                                                                                     
        global_tmr_voter(0)(118)  <=    (tmr_registers(0)(118) and tmr_registers(1)(118)) or                                            
                            (tmr_registers(1)(118) and tmr_registers(2)(118)) or                                                       
                            (tmr_registers(0)(118) and tmr_registers(2)(118));                                                         
                                                                                                                                     
        global_tmr_voter(0)(119)  <=    (tmr_registers(0)(119) and tmr_registers(1)(119)) or                                            
                            (tmr_registers(1)(119) and tmr_registers(2)(119)) or                                                       
                            (tmr_registers(0)(119) and tmr_registers(2)(119));                                                         
                                                                                                                                     
        global_tmr_voter(0)(120)  <=    (tmr_registers(0)(120) and tmr_registers(1)(120)) or                                            
                            (tmr_registers(1)(120) and tmr_registers(2)(120)) or                                                       
                            (tmr_registers(0)(120) and tmr_registers(2)(120));                                                         
                                                                                                                                     
        global_tmr_voter(0)(121)  <=    (tmr_registers(0)(121) and tmr_registers(1)(121)) or                                            
                            (tmr_registers(1)(121) and tmr_registers(2)(121)) or                                                       
                            (tmr_registers(0)(121) and tmr_registers(2)(121));                                                         
                                                                                                                                     
        global_tmr_voter(0)(122)  <=    (tmr_registers(0)(122) and tmr_registers(1)(122)) or                                            
                            (tmr_registers(1)(122) and tmr_registers(2)(122)) or                                                       
                            (tmr_registers(0)(122) and tmr_registers(2)(122));                                                         
                                                                                                                                     
        global_tmr_voter(0)(123)  <=    (tmr_registers(0)(123) and tmr_registers(1)(123)) or                                            
                            (tmr_registers(1)(123) and tmr_registers(2)(123)) or                                                       
                            (tmr_registers(0)(123) and tmr_registers(2)(123));                                                         
                                                                                                                                     
        global_tmr_voter(0)(124)  <=    (tmr_registers(0)(124) and tmr_registers(1)(124)) or                                            
                            (tmr_registers(1)(124) and tmr_registers(2)(124)) or                                                       
                            (tmr_registers(0)(124) and tmr_registers(2)(124));                                                         
                                                                                                                                     
        global_tmr_voter(0)(125)  <=    (tmr_registers(0)(125) and tmr_registers(1)(125)) or                                            
                            (tmr_registers(1)(125) and tmr_registers(2)(125)) or                                                       
                            (tmr_registers(0)(125) and tmr_registers(2)(125));                                                         
                                                                                                                                     
        global_tmr_voter(0)(126)  <=    (tmr_registers(0)(126) and tmr_registers(1)(126)) or                                            
                            (tmr_registers(1)(126) and tmr_registers(2)(126)) or                                                       
                            (tmr_registers(0)(126) and tmr_registers(2)(126));                                                         
                                                                                                                                     
        global_tmr_voter(0)(127)  <=    (tmr_registers(0)(127) and tmr_registers(1)(127)) or                                            
                            (tmr_registers(1)(127) and tmr_registers(2)(127)) or                                                       
                            (tmr_registers(0)(127) and tmr_registers(2)(127));                                                         
                                                                                                                                     
        global_tmr_voter(0)(128)  <=    (tmr_registers(0)(128) and tmr_registers(1)(128)) or                                            
                            (tmr_registers(1)(128) and tmr_registers(2)(128)) or                                                       
                            (tmr_registers(0)(128) and tmr_registers(2)(128));                                                         
                                                                                                                                     
        global_tmr_voter(0)(129)  <=    (tmr_registers(0)(129) and tmr_registers(1)(129)) or                                            
                            (tmr_registers(1)(129) and tmr_registers(2)(129)) or                                                       
                            (tmr_registers(0)(129) and tmr_registers(2)(129));                                                         
                                                                                                                                     
        global_tmr_voter(0)(130)  <=    (tmr_registers(0)(130) and tmr_registers(1)(130)) or                                            
                            (tmr_registers(1)(130) and tmr_registers(2)(130)) or                                                       
                            (tmr_registers(0)(130) and tmr_registers(2)(130));                                                         
                                                                                                                                     
        global_tmr_voter(0)(131)  <=    (tmr_registers(0)(131) and tmr_registers(1)(131)) or                                            
                            (tmr_registers(1)(131) and tmr_registers(2)(131)) or                                                       
                            (tmr_registers(0)(131) and tmr_registers(2)(131));                                                         
                                                                                                                                     
        global_tmr_voter(0)(132)  <=    (tmr_registers(0)(132) and tmr_registers(1)(132)) or                                            
                            (tmr_registers(1)(132) and tmr_registers(2)(132)) or                                                       
                            (tmr_registers(0)(132) and tmr_registers(2)(132));                                                         
                                                                                                                                     
        global_tmr_voter(0)(133)  <=    (tmr_registers(0)(133) and tmr_registers(1)(133)) or                                            
                            (tmr_registers(1)(133) and tmr_registers(2)(133)) or                                                       
                            (tmr_registers(0)(133) and tmr_registers(2)(133));                                                         
                                                                                                                                     
        global_tmr_voter(0)(134)  <=    (tmr_registers(0)(134) and tmr_registers(1)(134)) or                                            
                            (tmr_registers(1)(134) and tmr_registers(2)(134)) or                                                       
                            (tmr_registers(0)(134) and tmr_registers(2)(134));                                                         
                                                                                                                                     
        global_tmr_voter(0)(135)  <=    (tmr_registers(0)(135) and tmr_registers(1)(135)) or                                            
                            (tmr_registers(1)(135) and tmr_registers(2)(135)) or                                                       
                            (tmr_registers(0)(135) and tmr_registers(2)(135));                                                         
                                                                                                                                     
        global_tmr_voter(0)(136)  <=    (tmr_registers(0)(136) and tmr_registers(1)(136)) or                                            
                            (tmr_registers(1)(136) and tmr_registers(2)(136)) or                                                       
                            (tmr_registers(0)(136) and tmr_registers(2)(136));                                                         
                                                                                                                                     
        global_tmr_voter(0)(137)  <=    (tmr_registers(0)(137) and tmr_registers(1)(137)) or                                            
                            (tmr_registers(1)(137) and tmr_registers(2)(137)) or                                                       
                            (tmr_registers(0)(137) and tmr_registers(2)(137));                                                         
                                                                                                                                     
        global_tmr_voter(0)(138)  <=    (tmr_registers(0)(138) and tmr_registers(1)(138)) or                                            
                            (tmr_registers(1)(138) and tmr_registers(2)(138)) or                                                       
                            (tmr_registers(0)(138) and tmr_registers(2)(138));                                                         
                                                                                                                                     
        global_tmr_voter(0)(139)  <=    (tmr_registers(0)(139) and tmr_registers(1)(139)) or                                            
                            (tmr_registers(1)(139) and tmr_registers(2)(139)) or                                                       
                            (tmr_registers(0)(139) and tmr_registers(2)(139));                                                         
                                                                                                                                     
        global_tmr_voter(0)(140)  <=    (tmr_registers(0)(140) and tmr_registers(1)(140)) or                                            
                            (tmr_registers(1)(140) and tmr_registers(2)(140)) or                                                       
                            (tmr_registers(0)(140) and tmr_registers(2)(140));                                                         
                                                                                                                                     
        global_tmr_voter(0)(141)  <=    (tmr_registers(0)(141) and tmr_registers(1)(141)) or                                            
                            (tmr_registers(1)(141) and tmr_registers(2)(141)) or                                                       
                            (tmr_registers(0)(141) and tmr_registers(2)(141));                                                         
                                                                                                                                     
        global_tmr_voter(0)(142)  <=    (tmr_registers(0)(142) and tmr_registers(1)(142)) or                                            
                            (tmr_registers(1)(142) and tmr_registers(2)(142)) or                                                       
                            (tmr_registers(0)(142) and tmr_registers(2)(142));                                                         
                                                                                                                                     
        global_tmr_voter(0)(143)  <=    (tmr_registers(0)(143) and tmr_registers(1)(143)) or                                            
                            (tmr_registers(1)(143) and tmr_registers(2)(143)) or                                                       
                            (tmr_registers(0)(143) and tmr_registers(2)(143));                                                         
                                                                                                                                     
        global_tmr_voter(0)(144)  <=    (tmr_registers(0)(144) and tmr_registers(1)(144)) or                                            
                            (tmr_registers(1)(144) and tmr_registers(2)(144)) or                                                       
                            (tmr_registers(0)(144) and tmr_registers(2)(144));                                                         
                                                                                                                                     
        global_tmr_voter(0)(145)  <=    (tmr_registers(0)(145) and tmr_registers(1)(145)) or                                            
                            (tmr_registers(1)(145) and tmr_registers(2)(145)) or                                                       
                            (tmr_registers(0)(145) and tmr_registers(2)(145));                                                         
                                                                                                                                     
        global_tmr_voter(0)(146)  <=    (tmr_registers(0)(146) and tmr_registers(1)(146)) or                                            
                            (tmr_registers(1)(146) and tmr_registers(2)(146)) or                                                       
                            (tmr_registers(0)(146) and tmr_registers(2)(146));                                                         
                                                                                                                                     
        global_tmr_voter(0)(147)  <=    (tmr_registers(0)(147) and tmr_registers(1)(147)) or                                            
                            (tmr_registers(1)(147) and tmr_registers(2)(147)) or                                                       
                            (tmr_registers(0)(147) and tmr_registers(2)(147));                                                         
                                                                                                                                     
        global_tmr_voter(0)(148)  <=    (tmr_registers(0)(148) and tmr_registers(1)(148)) or                                            
                            (tmr_registers(1)(148) and tmr_registers(2)(148)) or                                                       
                            (tmr_registers(0)(148) and tmr_registers(2)(148));                                                         
                                                                                                                                     
        global_tmr_voter(0)(149)  <=    (tmr_registers(0)(149) and tmr_registers(1)(149)) or                                            
                            (tmr_registers(1)(149) and tmr_registers(2)(149)) or                                                       
                            (tmr_registers(0)(149) and tmr_registers(2)(149));                                                         
                                                                                                                                     
        global_tmr_voter(0)(150)  <=    (tmr_registers(0)(150) and tmr_registers(1)(150)) or                                            
                            (tmr_registers(1)(150) and tmr_registers(2)(150)) or                                                       
                            (tmr_registers(0)(150) and tmr_registers(2)(150));                                                         
                                                                                                                                     
        global_tmr_voter(0)(151)  <=    (tmr_registers(0)(151) and tmr_registers(1)(151)) or                                            
                            (tmr_registers(1)(151) and tmr_registers(2)(151)) or                                                       
                            (tmr_registers(0)(151) and tmr_registers(2)(151));                                                         
                                                                                                                                     
        global_tmr_voter(0)(152)  <=    (tmr_registers(0)(152) and tmr_registers(1)(152)) or                                            
                            (tmr_registers(1)(152) and tmr_registers(2)(152)) or                                                       
                            (tmr_registers(0)(152) and tmr_registers(2)(152));                                                         
                                                                                                                                     
        global_tmr_voter(0)(153)  <=    (tmr_registers(0)(153) and tmr_registers(1)(153)) or                                            
                            (tmr_registers(1)(153) and tmr_registers(2)(153)) or                                                       
                            (tmr_registers(0)(153) and tmr_registers(2)(153));                                                         
                                                                                                                                     
        global_tmr_voter(0)(154)  <=    (tmr_registers(0)(154) and tmr_registers(1)(154)) or                                            
                            (tmr_registers(1)(154) and tmr_registers(2)(154)) or                                                       
                            (tmr_registers(0)(154) and tmr_registers(2)(154));                                                         
                                                                                                                                     
        global_tmr_voter(0)(155)  <=    (tmr_registers(0)(155) and tmr_registers(1)(155)) or                                            
                            (tmr_registers(1)(155) and tmr_registers(2)(155)) or                                                       
                            (tmr_registers(0)(155) and tmr_registers(2)(155));                                                         
                                                                                                                                     
        global_tmr_voter(0)(156)  <=    (tmr_registers(0)(156) and tmr_registers(1)(156)) or                                            
                            (tmr_registers(1)(156) and tmr_registers(2)(156)) or                                                       
                            (tmr_registers(0)(156) and tmr_registers(2)(156));                                                         
                                                                                                                                     
        global_tmr_voter(0)(157)  <=    (tmr_registers(0)(157) and tmr_registers(1)(157)) or                                            
                            (tmr_registers(1)(157) and tmr_registers(2)(157)) or                                                       
                            (tmr_registers(0)(157) and tmr_registers(2)(157));                                                         
                                                                                                                                     
        global_tmr_voter(0)(158)  <=    (tmr_registers(0)(158) and tmr_registers(1)(158)) or                                            
                            (tmr_registers(1)(158) and tmr_registers(2)(158)) or                                                       
                            (tmr_registers(0)(158) and tmr_registers(2)(158));                                                         
                                                                                                                                     
        global_tmr_voter(0)(159)  <=    (tmr_registers(0)(159) and tmr_registers(1)(159)) or                                            
                            (tmr_registers(1)(159) and tmr_registers(2)(159)) or                                                       
                            (tmr_registers(0)(159) and tmr_registers(2)(159));                                                         
                                                                                                                                     
        global_tmr_voter(0)(160)  <=    (tmr_registers(0)(160) and tmr_registers(1)(160)) or                                            
                            (tmr_registers(1)(160) and tmr_registers(2)(160)) or                                                       
                            (tmr_registers(0)(160) and tmr_registers(2)(160));                                                         
                                                                                                                                     
        global_tmr_voter(0)(161)  <=    (tmr_registers(0)(161) and tmr_registers(1)(161)) or                                            
                            (tmr_registers(1)(161) and tmr_registers(2)(161)) or                                                       
                            (tmr_registers(0)(161) and tmr_registers(2)(161));                                                         
                                                                                                                                     
        global_tmr_voter(0)(162)  <=    (tmr_registers(0)(162) and tmr_registers(1)(162)) or                                            
                            (tmr_registers(1)(162) and tmr_registers(2)(162)) or                                                       
                            (tmr_registers(0)(162) and tmr_registers(2)(162));                                                         
                                                                                                                                     
        global_tmr_voter(0)(163)  <=    (tmr_registers(0)(163) and tmr_registers(1)(163)) or                                            
                            (tmr_registers(1)(163) and tmr_registers(2)(163)) or                                                       
                            (tmr_registers(0)(163) and tmr_registers(2)(163));                                                         
                                                                                                                                     
        global_tmr_voter(0)(164)  <=    (tmr_registers(0)(164) and tmr_registers(1)(164)) or                                            
                            (tmr_registers(1)(164) and tmr_registers(2)(164)) or                                                       
                            (tmr_registers(0)(164) and tmr_registers(2)(164));                                                         
                                                                                                                                     
        global_tmr_voter(0)(165)  <=    (tmr_registers(0)(165) and tmr_registers(1)(165)) or                                            
                            (tmr_registers(1)(165) and tmr_registers(2)(165)) or                                                       
                            (tmr_registers(0)(165) and tmr_registers(2)(165));                                                         
                                                                                                                                     
        global_tmr_voter(0)(166)  <=    (tmr_registers(0)(166) and tmr_registers(1)(166)) or                                            
                            (tmr_registers(1)(166) and tmr_registers(2)(166)) or                                                       
                            (tmr_registers(0)(166) and tmr_registers(2)(166));                                                         
                                                                                                                                     
        global_tmr_voter(0)(167)  <=    (tmr_registers(0)(167) and tmr_registers(1)(167)) or                                            
                            (tmr_registers(1)(167) and tmr_registers(2)(167)) or                                                       
                            (tmr_registers(0)(167) and tmr_registers(2)(167));                                                         
                                                                                                                                     
        global_tmr_voter(0)(168)  <=    (tmr_registers(0)(168) and tmr_registers(1)(168)) or                                            
                            (tmr_registers(1)(168) and tmr_registers(2)(168)) or                                                       
                            (tmr_registers(0)(168) and tmr_registers(2)(168));                                                         
                                                                                                                                     
        global_tmr_voter(0)(169)  <=    (tmr_registers(0)(169) and tmr_registers(1)(169)) or                                            
                            (tmr_registers(1)(169) and tmr_registers(2)(169)) or                                                       
                            (tmr_registers(0)(169) and tmr_registers(2)(169));                                                         
                                                                                                                                     
        global_tmr_voter(0)(170)  <=    (tmr_registers(0)(170) and tmr_registers(1)(170)) or                                            
                            (tmr_registers(1)(170) and tmr_registers(2)(170)) or                                                       
                            (tmr_registers(0)(170) and tmr_registers(2)(170));                                                         
                                                                                                                                     
        global_tmr_voter(0)(171)  <=    (tmr_registers(0)(171) and tmr_registers(1)(171)) or                                            
                            (tmr_registers(1)(171) and tmr_registers(2)(171)) or                                                       
                            (tmr_registers(0)(171) and tmr_registers(2)(171));                                                         
                                                                                                                                     
        global_tmr_voter(0)(172)  <=    (tmr_registers(0)(172) and tmr_registers(1)(172)) or                                            
                            (tmr_registers(1)(172) and tmr_registers(2)(172)) or                                                       
                            (tmr_registers(0)(172) and tmr_registers(2)(172));                                                         
                                                                                                                                     
        global_tmr_voter(0)(173)  <=    (tmr_registers(0)(173) and tmr_registers(1)(173)) or                                            
                            (tmr_registers(1)(173) and tmr_registers(2)(173)) or                                                       
                            (tmr_registers(0)(173) and tmr_registers(2)(173));                                                         
                                                                                                                                     
        global_tmr_voter(0)(174)  <=    (tmr_registers(0)(174) and tmr_registers(1)(174)) or                                            
                            (tmr_registers(1)(174) and tmr_registers(2)(174)) or                                                       
                            (tmr_registers(0)(174) and tmr_registers(2)(174));                                                         
                                                                                                                                     
        global_tmr_voter(0)(175)  <=    (tmr_registers(0)(175) and tmr_registers(1)(175)) or                                            
                            (tmr_registers(1)(175) and tmr_registers(2)(175)) or                                                       
                            (tmr_registers(0)(175) and tmr_registers(2)(175));                                                         
                                                                                                                                     
        global_tmr_voter(0)(176)  <=    (tmr_registers(0)(176) and tmr_registers(1)(176)) or                                            
                            (tmr_registers(1)(176) and tmr_registers(2)(176)) or                                                       
                            (tmr_registers(0)(176) and tmr_registers(2)(176));                                                         
                                                                                                                                     
        global_tmr_voter(0)(177)  <=    (tmr_registers(0)(177) and tmr_registers(1)(177)) or                                            
                            (tmr_registers(1)(177) and tmr_registers(2)(177)) or                                                       
                            (tmr_registers(0)(177) and tmr_registers(2)(177));                                                         
                                                                                                                                     
        global_tmr_voter(0)(178)  <=    (tmr_registers(0)(178) and tmr_registers(1)(178)) or                                            
                            (tmr_registers(1)(178) and tmr_registers(2)(178)) or                                                       
                            (tmr_registers(0)(178) and tmr_registers(2)(178));                                                         
                                                                                                                                     
        global_tmr_voter(0)(179)  <=    (tmr_registers(0)(179) and tmr_registers(1)(179)) or                                            
                            (tmr_registers(1)(179) and tmr_registers(2)(179)) or                                                       
                            (tmr_registers(0)(179) and tmr_registers(2)(179));                                                         
                                                                                                                                     
        global_tmr_voter(0)(180)  <=    (tmr_registers(0)(180) and tmr_registers(1)(180)) or                                            
                            (tmr_registers(1)(180) and tmr_registers(2)(180)) or                                                       
                            (tmr_registers(0)(180) and tmr_registers(2)(180));                                                         
                                                                                                                                     
        global_tmr_voter(0)(181)  <=    (tmr_registers(0)(181) and tmr_registers(1)(181)) or                                            
                            (tmr_registers(1)(181) and tmr_registers(2)(181)) or                                                       
                            (tmr_registers(0)(181) and tmr_registers(2)(181));                                                         
                                                                                                                                     
        global_tmr_voter(0)(182)  <=    (tmr_registers(0)(182) and tmr_registers(1)(182)) or                                            
                            (tmr_registers(1)(182) and tmr_registers(2)(182)) or                                                       
                            (tmr_registers(0)(182) and tmr_registers(2)(182));                                                         
                                                                                                                                     
        global_tmr_voter(0)(183)  <=    (tmr_registers(0)(183) and tmr_registers(1)(183)) or                                            
                            (tmr_registers(1)(183) and tmr_registers(2)(183)) or                                                       
                            (tmr_registers(0)(183) and tmr_registers(2)(183));                                                         
                                                                                                                                     
        global_tmr_voter(0)(184)  <=    (tmr_registers(0)(184) and tmr_registers(1)(184)) or                                            
                            (tmr_registers(1)(184) and tmr_registers(2)(184)) or                                                       
                            (tmr_registers(0)(184) and tmr_registers(2)(184));                                                         
                                                                                                                                     
        global_tmr_voter(0)(185)  <=    (tmr_registers(0)(185) and tmr_registers(1)(185)) or                                            
                            (tmr_registers(1)(185) and tmr_registers(2)(185)) or                                                       
                            (tmr_registers(0)(185) and tmr_registers(2)(185));                                                         
                                                                                                                                     
        global_tmr_voter(0)(186)  <=    (tmr_registers(0)(186) and tmr_registers(1)(186)) or                                            
                            (tmr_registers(1)(186) and tmr_registers(2)(186)) or                                                       
                            (tmr_registers(0)(186) and tmr_registers(2)(186));                                                         
                                                                                                                                     
        global_tmr_voter(0)(187)  <=    (tmr_registers(0)(187) and tmr_registers(1)(187)) or                                            
                            (tmr_registers(1)(187) and tmr_registers(2)(187)) or                                                       
                            (tmr_registers(0)(187) and tmr_registers(2)(187));                                                         
                                                                                                                                     
        global_tmr_voter(0)(188)  <=    (tmr_registers(0)(188) and tmr_registers(1)(188)) or                                            
                            (tmr_registers(1)(188) and tmr_registers(2)(188)) or                                                       
                            (tmr_registers(0)(188) and tmr_registers(2)(188));                                                         
                                                                                                                                     
        global_tmr_voter(0)(189)  <=    (tmr_registers(0)(189) and tmr_registers(1)(189)) or                                            
                            (tmr_registers(1)(189) and tmr_registers(2)(189)) or                                                       
                            (tmr_registers(0)(189) and tmr_registers(2)(189));                                                         
                                                                                                                                     
        global_tmr_voter(0)(190)  <=    (tmr_registers(0)(190) and tmr_registers(1)(190)) or                                            
                            (tmr_registers(1)(190) and tmr_registers(2)(190)) or                                                       
                            (tmr_registers(0)(190) and tmr_registers(2)(190));                                                         
                                                                                                                                     
        global_tmr_voter(0)(191)  <=    (tmr_registers(0)(191) and tmr_registers(1)(191)) or                                            
                            (tmr_registers(1)(191) and tmr_registers(2)(191)) or                                                       
                            (tmr_registers(0)(191) and tmr_registers(2)(191));                                                         
                                                                                                                                     
        global_tmr_voter(0)(192)  <=    (tmr_registers(0)(192) and tmr_registers(1)(192)) or                                            
                            (tmr_registers(1)(192) and tmr_registers(2)(192)) or                                                       
                            (tmr_registers(0)(192) and tmr_registers(2)(192));                                                         
                                                                                                                                     
        global_tmr_voter(0)(193)  <=    (tmr_registers(0)(193) and tmr_registers(1)(193)) or                                            
                            (tmr_registers(1)(193) and tmr_registers(2)(193)) or                                                       
                            (tmr_registers(0)(193) and tmr_registers(2)(193));                                                         
                                                                                                                                     
        global_tmr_voter(0)(194)  <=    (tmr_registers(0)(194) and tmr_registers(1)(194)) or                                            
                            (tmr_registers(1)(194) and tmr_registers(2)(194)) or                                                       
                            (tmr_registers(0)(194) and tmr_registers(2)(194));                                                         
                                                                                                                                     
        global_tmr_voter(0)(195)  <=    (tmr_registers(0)(195) and tmr_registers(1)(195)) or                                            
                            (tmr_registers(1)(195) and tmr_registers(2)(195)) or                                                       
                            (tmr_registers(0)(195) and tmr_registers(2)(195));                                                         
                                                                                                                                     
        global_tmr_voter(0)(196)  <=    (tmr_registers(0)(196) and tmr_registers(1)(196)) or                                            
                            (tmr_registers(1)(196) and tmr_registers(2)(196)) or                                                       
                            (tmr_registers(0)(196) and tmr_registers(2)(196));                                                         
                                                                                                                                     
        global_tmr_voter(0)(197)  <=    (tmr_registers(0)(197) and tmr_registers(1)(197)) or                                            
                            (tmr_registers(1)(197) and tmr_registers(2)(197)) or                                                       
                            (tmr_registers(0)(197) and tmr_registers(2)(197));                                                         
                                                                                                                                     
        global_tmr_voter(0)(198)  <=    (tmr_registers(0)(198) and tmr_registers(1)(198)) or                                            
                            (tmr_registers(1)(198) and tmr_registers(2)(198)) or                                                       
                            (tmr_registers(0)(198) and tmr_registers(2)(198));                                                         
                                                                                                                                     
        global_tmr_voter(0)(199)  <=    (tmr_registers(0)(199) and tmr_registers(1)(199)) or                                            
                            (tmr_registers(1)(199) and tmr_registers(2)(199)) or                                                       
                            (tmr_registers(0)(199) and tmr_registers(2)(199));                                                         
                                                                                                                                     
        global_tmr_voter(0)(200)  <=    (tmr_registers(0)(200) and tmr_registers(1)(200)) or                                            
                            (tmr_registers(1)(200) and tmr_registers(2)(200)) or                                                       
                            (tmr_registers(0)(200) and tmr_registers(2)(200));                                                         
                                                                                                                                     
        global_tmr_voter(0)(201)  <=    (tmr_registers(0)(201) and tmr_registers(1)(201)) or                                            
                            (tmr_registers(1)(201) and tmr_registers(2)(201)) or                                                       
                            (tmr_registers(0)(201) and tmr_registers(2)(201));                                                         
                                                                                                                                     
        global_tmr_voter(0)(202)  <=    (tmr_registers(0)(202) and tmr_registers(1)(202)) or                                            
                            (tmr_registers(1)(202) and tmr_registers(2)(202)) or                                                       
                            (tmr_registers(0)(202) and tmr_registers(2)(202));                                                         
                                                                                                                                     
        global_tmr_voter(0)(203)  <=    (tmr_registers(0)(203) and tmr_registers(1)(203)) or                                            
                            (tmr_registers(1)(203) and tmr_registers(2)(203)) or                                                       
                            (tmr_registers(0)(203) and tmr_registers(2)(203));                                                         
                                                                                                                                     
        global_tmr_voter(0)(204)  <=    (tmr_registers(0)(204) and tmr_registers(1)(204)) or                                            
                            (tmr_registers(1)(204) and tmr_registers(2)(204)) or                                                       
                            (tmr_registers(0)(204) and tmr_registers(2)(204));                                                         
                                                                                                                                     
        global_tmr_voter(0)(205)  <=    (tmr_registers(0)(205) and tmr_registers(1)(205)) or                                            
                            (tmr_registers(1)(205) and tmr_registers(2)(205)) or                                                       
                            (tmr_registers(0)(205) and tmr_registers(2)(205));                                                         
                                                                                                                                     
        global_tmr_voter(0)(206)  <=    (tmr_registers(0)(206) and tmr_registers(1)(206)) or                                            
                            (tmr_registers(1)(206) and tmr_registers(2)(206)) or                                                       
                            (tmr_registers(0)(206) and tmr_registers(2)(206));                                                         
                                                                                                                                     
        global_tmr_voter(0)(207)  <=    (tmr_registers(0)(207) and tmr_registers(1)(207)) or                                            
                            (tmr_registers(1)(207) and tmr_registers(2)(207)) or                                                       
                            (tmr_registers(0)(207) and tmr_registers(2)(207));                                                         
                                                                                                                                     
        global_tmr_voter(0)(208)  <=    (tmr_registers(0)(208) and tmr_registers(1)(208)) or                                            
                            (tmr_registers(1)(208) and tmr_registers(2)(208)) or                                                       
                            (tmr_registers(0)(208) and tmr_registers(2)(208));                                                         
                                                                                                                                     
        global_tmr_voter(0)(209)  <=    (tmr_registers(0)(209) and tmr_registers(1)(209)) or                                            
                            (tmr_registers(1)(209) and tmr_registers(2)(209)) or                                                       
                            (tmr_registers(0)(209) and tmr_registers(2)(209));                                                         
                                                                                                                                     
        global_tmr_voter(0)(210)  <=    (tmr_registers(0)(210) and tmr_registers(1)(210)) or                                            
                            (tmr_registers(1)(210) and tmr_registers(2)(210)) or                                                       
                            (tmr_registers(0)(210) and tmr_registers(2)(210));                                                         
                                                                                                                                     
        global_tmr_voter(0)(211)  <=    (tmr_registers(0)(211) and tmr_registers(1)(211)) or                                            
                            (tmr_registers(1)(211) and tmr_registers(2)(211)) or                                                       
                            (tmr_registers(0)(211) and tmr_registers(2)(211));                                                         
                                                                                                                                     
        global_tmr_voter(0)(212)  <=    (tmr_registers(0)(212) and tmr_registers(1)(212)) or                                            
                            (tmr_registers(1)(212) and tmr_registers(2)(212)) or                                                       
                            (tmr_registers(0)(212) and tmr_registers(2)(212));                                                         
                                                                                                                                     
        global_tmr_voter(0)(213)  <=    (tmr_registers(0)(213) and tmr_registers(1)(213)) or                                            
                            (tmr_registers(1)(213) and tmr_registers(2)(213)) or                                                       
                            (tmr_registers(0)(213) and tmr_registers(2)(213));                                                         
                                                                                                                                     
        global_tmr_voter(0)(214)  <=    (tmr_registers(0)(214) and tmr_registers(1)(214)) or                                            
                            (tmr_registers(1)(214) and tmr_registers(2)(214)) or                                                       
                            (tmr_registers(0)(214) and tmr_registers(2)(214));                                                         
                                                                                                                                     
        global_tmr_voter(0)(215)  <=    (tmr_registers(0)(215) and tmr_registers(1)(215)) or                                            
                            (tmr_registers(1)(215) and tmr_registers(2)(215)) or                                                       
                            (tmr_registers(0)(215) and tmr_registers(2)(215));                                                         
                                                                                                                                     
        global_tmr_voter(0)(216)  <=    (tmr_registers(0)(216) and tmr_registers(1)(216)) or                                            
                            (tmr_registers(1)(216) and tmr_registers(2)(216)) or                                                       
                            (tmr_registers(0)(216) and tmr_registers(2)(216));                                                         
                                                                                                                                     
        global_tmr_voter(0)(217)  <=    (tmr_registers(0)(217) and tmr_registers(1)(217)) or                                            
                            (tmr_registers(1)(217) and tmr_registers(2)(217)) or                                                       
                            (tmr_registers(0)(217) and tmr_registers(2)(217));                                                         
                                                                                                                                     
        global_tmr_voter(0)(218)  <=    (tmr_registers(0)(218) and tmr_registers(1)(218)) or                                            
                            (tmr_registers(1)(218) and tmr_registers(2)(218)) or                                                       
                            (tmr_registers(0)(218) and tmr_registers(2)(218));                                                         
                                                                                                                                     
        global_tmr_voter(0)(219)  <=    (tmr_registers(0)(219) and tmr_registers(1)(219)) or                                            
                            (tmr_registers(1)(219) and tmr_registers(2)(219)) or                                                       
                            (tmr_registers(0)(219) and tmr_registers(2)(219));                                                         
                                                                                                                                     
        global_tmr_voter(0)(220)  <=    (tmr_registers(0)(220) and tmr_registers(1)(220)) or                                            
                            (tmr_registers(1)(220) and tmr_registers(2)(220)) or                                                       
                            (tmr_registers(0)(220) and tmr_registers(2)(220));                                                         
                                                                                                                                     
        global_tmr_voter(0)(221)  <=    (tmr_registers(0)(221) and tmr_registers(1)(221)) or                                            
                            (tmr_registers(1)(221) and tmr_registers(2)(221)) or                                                       
                            (tmr_registers(0)(221) and tmr_registers(2)(221));                                                         
                                                                                                                                     
        global_tmr_voter(0)(222)  <=    (tmr_registers(0)(222) and tmr_registers(1)(222)) or                                            
                            (tmr_registers(1)(222) and tmr_registers(2)(222)) or                                                       
                            (tmr_registers(0)(222) and tmr_registers(2)(222));                                                         
                                                                                                                                     
        global_tmr_voter(0)(223)  <=    (tmr_registers(0)(223) and tmr_registers(1)(223)) or                                            
                            (tmr_registers(1)(223) and tmr_registers(2)(223)) or                                                       
                            (tmr_registers(0)(223) and tmr_registers(2)(223));                                                         
                                                                                                                                     
        global_tmr_voter(0)(224)  <=    (tmr_registers(0)(224) and tmr_registers(1)(224)) or                                            
                            (tmr_registers(1)(224) and tmr_registers(2)(224)) or                                                       
                            (tmr_registers(0)(224) and tmr_registers(2)(224));                                                         
                                                                                                                                     
        global_tmr_voter(0)(225)  <=    (tmr_registers(0)(225) and tmr_registers(1)(225)) or                                            
                            (tmr_registers(1)(225) and tmr_registers(2)(225)) or                                                       
                            (tmr_registers(0)(225) and tmr_registers(2)(225));                                                         
                                                                                                                                     
        global_tmr_voter(0)(226)  <=    (tmr_registers(0)(226) and tmr_registers(1)(226)) or                                            
                            (tmr_registers(1)(226) and tmr_registers(2)(226)) or                                                       
                            (tmr_registers(0)(226) and tmr_registers(2)(226));                                                         
                                                                                                                                     
        global_tmr_voter(0)(227)  <=    (tmr_registers(0)(227) and tmr_registers(1)(227)) or                                            
                            (tmr_registers(1)(227) and tmr_registers(2)(227)) or                                                       
                            (tmr_registers(0)(227) and tmr_registers(2)(227));                                                         
                                                                                                                                     
        global_tmr_voter(0)(228)  <=    (tmr_registers(0)(228) and tmr_registers(1)(228)) or                                            
                            (tmr_registers(1)(228) and tmr_registers(2)(228)) or                                                       
                            (tmr_registers(0)(228) and tmr_registers(2)(228));                                                         
                                                                                                                                     
        global_tmr_voter(0)(229)  <=    (tmr_registers(0)(229) and tmr_registers(1)(229)) or                                            
                            (tmr_registers(1)(229) and tmr_registers(2)(229)) or                                                       
                            (tmr_registers(0)(229) and tmr_registers(2)(229));                                                         
                                                                                                                                     
        global_tmr_voter(0)(230)  <=    (tmr_registers(0)(230) and tmr_registers(1)(230)) or                                            
                            (tmr_registers(1)(230) and tmr_registers(2)(230)) or                                                       
                            (tmr_registers(0)(230) and tmr_registers(2)(230));                                                         
                                                                                                                                     
        global_tmr_voter(0)(231)  <=    (tmr_registers(0)(231) and tmr_registers(1)(231)) or                                            
                            (tmr_registers(1)(231) and tmr_registers(2)(231)) or                                                       
                            (tmr_registers(0)(231) and tmr_registers(2)(231));                                                         
                                                                                                                                     
        global_tmr_voter(0)(232)  <=    (tmr_registers(0)(232) and tmr_registers(1)(232)) or                                            
                            (tmr_registers(1)(232) and tmr_registers(2)(232)) or                                                       
                            (tmr_registers(0)(232) and tmr_registers(2)(232));                                                         
                                                                                                                                     
        global_tmr_voter(0)(233)  <=    (tmr_registers(0)(233) and tmr_registers(1)(233)) or                                            
                            (tmr_registers(1)(233) and tmr_registers(2)(233)) or                                                       
                            (tmr_registers(0)(233) and tmr_registers(2)(233));                                                         
                                                                                                                                     
        global_tmr_voter(0)(234)  <=    (tmr_registers(0)(234) and tmr_registers(1)(234)) or                                            
                            (tmr_registers(1)(234) and tmr_registers(2)(234)) or                                                       
                            (tmr_registers(0)(234) and tmr_registers(2)(234));                                                         
                                                                                                                                     
        global_tmr_voter(0)(235)  <=    (tmr_registers(0)(235) and tmr_registers(1)(235)) or                                            
                            (tmr_registers(1)(235) and tmr_registers(2)(235)) or                                                       
                            (tmr_registers(0)(235) and tmr_registers(2)(235));                                                         
                                                                                                                                     
        global_tmr_voter(0)(236)  <=    (tmr_registers(0)(236) and tmr_registers(1)(236)) or                                            
                            (tmr_registers(1)(236) and tmr_registers(2)(236)) or                                                       
                            (tmr_registers(0)(236) and tmr_registers(2)(236));                                                         
                                                                                                                                     
        global_tmr_voter(0)(237)  <=    (tmr_registers(0)(237) and tmr_registers(1)(237)) or                                            
                            (tmr_registers(1)(237) and tmr_registers(2)(237)) or                                                       
                            (tmr_registers(0)(237) and tmr_registers(2)(237));                                                         
                                                                                                                                     
        global_tmr_voter(0)(238)  <=    (tmr_registers(0)(238) and tmr_registers(1)(238)) or                                            
                            (tmr_registers(1)(238) and tmr_registers(2)(238)) or                                                       
                            (tmr_registers(0)(238) and tmr_registers(2)(238));                                                         
                                                                                                                                     
        global_tmr_voter(0)(239)  <=    (tmr_registers(0)(239) and tmr_registers(1)(239)) or                                            
                            (tmr_registers(1)(239) and tmr_registers(2)(239)) or                                                       
                            (tmr_registers(0)(239) and tmr_registers(2)(239));                                                         
                                                                                                                                     
        global_tmr_voter(0)(240)  <=    (tmr_registers(0)(240) and tmr_registers(1)(240)) or                                            
                            (tmr_registers(1)(240) and tmr_registers(2)(240)) or                                                       
                            (tmr_registers(0)(240) and tmr_registers(2)(240));                                                         
                                                                                                                                     
        global_tmr_voter(0)(241)  <=    (tmr_registers(0)(241) and tmr_registers(1)(241)) or                                            
                            (tmr_registers(1)(241) and tmr_registers(2)(241)) or                                                       
                            (tmr_registers(0)(241) and tmr_registers(2)(241));                                                         
                                                                                                                                     
        global_tmr_voter(0)(242)  <=    (tmr_registers(0)(242) and tmr_registers(1)(242)) or                                            
                            (tmr_registers(1)(242) and tmr_registers(2)(242)) or                                                       
                            (tmr_registers(0)(242) and tmr_registers(2)(242));                                                         
                                                                                                                                     
        global_tmr_voter(0)(243)  <=    (tmr_registers(0)(243) and tmr_registers(1)(243)) or                                            
                            (tmr_registers(1)(243) and tmr_registers(2)(243)) or                                                       
                            (tmr_registers(0)(243) and tmr_registers(2)(243));                                                         
                                                                                                                                     
        global_tmr_voter(0)(244)  <=    (tmr_registers(0)(244) and tmr_registers(1)(244)) or                                            
                            (tmr_registers(1)(244) and tmr_registers(2)(244)) or                                                       
                            (tmr_registers(0)(244) and tmr_registers(2)(244));                                                         
                                                                                                                                     
        global_tmr_voter(0)(245)  <=    (tmr_registers(0)(245) and tmr_registers(1)(245)) or                                            
                            (tmr_registers(1)(245) and tmr_registers(2)(245)) or                                                       
                            (tmr_registers(0)(245) and tmr_registers(2)(245));                                                         
                                                                                                                                     
        global_tmr_voter(0)(246)  <=    (tmr_registers(0)(246) and tmr_registers(1)(246)) or                                            
                            (tmr_registers(1)(246) and tmr_registers(2)(246)) or                                                       
                            (tmr_registers(0)(246) and tmr_registers(2)(246));                                                         
                                                                                                                                     
        global_tmr_voter(0)(247)  <=    (tmr_registers(0)(247) and tmr_registers(1)(247)) or                                            
                            (tmr_registers(1)(247) and tmr_registers(2)(247)) or                                                       
                            (tmr_registers(0)(247) and tmr_registers(2)(247));                                                         
                                                                                                                                     
        global_tmr_voter(0)(248)  <=    (tmr_registers(0)(248) and tmr_registers(1)(248)) or                                            
                            (tmr_registers(1)(248) and tmr_registers(2)(248)) or                                                       
                            (tmr_registers(0)(248) and tmr_registers(2)(248));                                                         
                                                                                                                                     
        global_tmr_voter(0)(249)  <=    (tmr_registers(0)(249) and tmr_registers(1)(249)) or                                            
                            (tmr_registers(1)(249) and tmr_registers(2)(249)) or                                                       
                            (tmr_registers(0)(249) and tmr_registers(2)(249));                                                         
                                                                                                                                     
        global_tmr_voter(0)(250)  <=    (tmr_registers(0)(250) and tmr_registers(1)(250)) or                                            
                            (tmr_registers(1)(250) and tmr_registers(2)(250)) or                                                       
                            (tmr_registers(0)(250) and tmr_registers(2)(250));                                                         
                                                                                                                                     
        global_tmr_voter(0)(251)  <=    (tmr_registers(0)(251) and tmr_registers(1)(251)) or                                            
                            (tmr_registers(1)(251) and tmr_registers(2)(251)) or                                                       
                            (tmr_registers(0)(251) and tmr_registers(2)(251));                                                         
                                                                                                                                     
        global_tmr_voter(0)(252)  <=    (tmr_registers(0)(252) and tmr_registers(1)(252)) or                                            
                            (tmr_registers(1)(252) and tmr_registers(2)(252)) or                                                       
                            (tmr_registers(0)(252) and tmr_registers(2)(252));                                                         
                                                                                                                                     
        global_tmr_voter(0)(253)  <=    (tmr_registers(0)(253) and tmr_registers(1)(253)) or                                            
                            (tmr_registers(1)(253) and tmr_registers(2)(253)) or                                                       
                            (tmr_registers(0)(253) and tmr_registers(2)(253));                                                         
                                                                                                                                     
        global_tmr_voter(0)(254)  <=    (tmr_registers(0)(254) and tmr_registers(1)(254)) or                                            
                            (tmr_registers(1)(254) and tmr_registers(2)(254)) or                                                       
                            (tmr_registers(0)(254) and tmr_registers(2)(254));                                                         
                                                                                                                                     
        global_tmr_voter(0)(255)  <=    (tmr_registers(0)(255) and tmr_registers(1)(255)) or                                            
                            (tmr_registers(1)(255) and tmr_registers(2)(255)) or                                                       
                            (tmr_registers(0)(255) and tmr_registers(2)(255));                                                         
                                                                                                                                     
        global_tmr_voter(0)(256)  <=    (tmr_registers(0)(256) and tmr_registers(1)(256)) or                                            
                            (tmr_registers(1)(256) and tmr_registers(2)(256)) or                                                       
                            (tmr_registers(0)(256) and tmr_registers(2)(256));                                                         
                                                                                                                                     
        global_tmr_voter(0)(257)  <=    (tmr_registers(0)(257) and tmr_registers(1)(257)) or                                            
                            (tmr_registers(1)(257) and tmr_registers(2)(257)) or                                                       
                            (tmr_registers(0)(257) and tmr_registers(2)(257));                                                         
                                                                                                                                     
        global_tmr_voter(0)(258)  <=    (tmr_registers(0)(258) and tmr_registers(1)(258)) or                                            
                            (tmr_registers(1)(258) and tmr_registers(2)(258)) or                                                       
                            (tmr_registers(0)(258) and tmr_registers(2)(258));                                                         
                                                                                                                                     
        global_tmr_voter(0)(259)  <=    (tmr_registers(0)(259) and tmr_registers(1)(259)) or                                            
                            (tmr_registers(1)(259) and tmr_registers(2)(259)) or                                                       
                            (tmr_registers(0)(259) and tmr_registers(2)(259));                                                         
                                                                                                                                     
        global_tmr_voter(0)(260)  <=    (tmr_registers(0)(260) and tmr_registers(1)(260)) or                                            
                            (tmr_registers(1)(260) and tmr_registers(2)(260)) or                                                       
                            (tmr_registers(0)(260) and tmr_registers(2)(260));                                                         
                                                                                                                                     
        global_tmr_voter(0)(261)  <=    (tmr_registers(0)(261) and tmr_registers(1)(261)) or                                            
                            (tmr_registers(1)(261) and tmr_registers(2)(261)) or                                                       
                            (tmr_registers(0)(261) and tmr_registers(2)(261));                                                         
                                                                                                                                     
        global_tmr_voter(0)(262)  <=    (tmr_registers(0)(262) and tmr_registers(1)(262)) or                                            
                            (tmr_registers(1)(262) and tmr_registers(2)(262)) or                                                       
                            (tmr_registers(0)(262) and tmr_registers(2)(262));                                                         
                                                                                                                                     
        global_tmr_voter(0)(263)  <=    (tmr_registers(0)(263) and tmr_registers(1)(263)) or                                            
                            (tmr_registers(1)(263) and tmr_registers(2)(263)) or                                                       
                            (tmr_registers(0)(263) and tmr_registers(2)(263));                                                         
                                                                                                                                     
        global_tmr_voter(0)(264)  <=    (tmr_registers(0)(264) and tmr_registers(1)(264)) or                                            
                            (tmr_registers(1)(264) and tmr_registers(2)(264)) or                                                       
                            (tmr_registers(0)(264) and tmr_registers(2)(264));                                                         
                                                                                                                                     
        global_tmr_voter(0)(265)  <=    (tmr_registers(0)(265) and tmr_registers(1)(265)) or                                            
                            (tmr_registers(1)(265) and tmr_registers(2)(265)) or                                                       
                            (tmr_registers(0)(265) and tmr_registers(2)(265));                                                         
                                                                                                                                     
        global_tmr_voter(0)(266)  <=    (tmr_registers(0)(266) and tmr_registers(1)(266)) or                                            
                            (tmr_registers(1)(266) and tmr_registers(2)(266)) or                                                       
                            (tmr_registers(0)(266) and tmr_registers(2)(266));                                                         
                                                                                                                                     
        global_tmr_voter(0)(267)  <=    (tmr_registers(0)(267) and tmr_registers(1)(267)) or                                            
                            (tmr_registers(1)(267) and tmr_registers(2)(267)) or                                                       
                            (tmr_registers(0)(267) and tmr_registers(2)(267));                                                         
                                                                                                                                     
        global_tmr_voter(0)(268)  <=    (tmr_registers(0)(268) and tmr_registers(1)(268)) or                                            
                            (tmr_registers(1)(268) and tmr_registers(2)(268)) or                                                       
                            (tmr_registers(0)(268) and tmr_registers(2)(268));                                                         
                                                                                                                                     
        global_tmr_voter(0)(269)  <=    (tmr_registers(0)(269) and tmr_registers(1)(269)) or                                            
                            (tmr_registers(1)(269) and tmr_registers(2)(269)) or                                                       
                            (tmr_registers(0)(269) and tmr_registers(2)(269));                                                         
                                                                                                                                     
        global_tmr_voter(0)(270)  <=    (tmr_registers(0)(270) and tmr_registers(1)(270)) or                                            
                            (tmr_registers(1)(270) and tmr_registers(2)(270)) or                                                       
                            (tmr_registers(0)(270) and tmr_registers(2)(270));                                                         
                                                                                                                                     
        global_tmr_voter(0)(271)  <=    (tmr_registers(0)(271) and tmr_registers(1)(271)) or                                            
                            (tmr_registers(1)(271) and tmr_registers(2)(271)) or                                                       
                            (tmr_registers(0)(271) and tmr_registers(2)(271));                                                         
                                                                                                                                     
        global_tmr_voter(0)(272)  <=    (tmr_registers(0)(272) and tmr_registers(1)(272)) or                                            
                            (tmr_registers(1)(272) and tmr_registers(2)(272)) or                                                       
                            (tmr_registers(0)(272) and tmr_registers(2)(272));                                                         
                                                                                                                                     
        global_tmr_voter(0)(273)  <=    (tmr_registers(0)(273) and tmr_registers(1)(273)) or                                            
                            (tmr_registers(1)(273) and tmr_registers(2)(273)) or                                                       
                            (tmr_registers(0)(273) and tmr_registers(2)(273));                                                         
                                                                                                                                     
        global_tmr_voter(0)(274)  <=    (tmr_registers(0)(274) and tmr_registers(1)(274)) or                                            
                            (tmr_registers(1)(274) and tmr_registers(2)(274)) or                                                       
                            (tmr_registers(0)(274) and tmr_registers(2)(274));                                                         
                                                                                                                                     
        global_tmr_voter(0)(275)  <=    (tmr_registers(0)(275) and tmr_registers(1)(275)) or                                            
                            (tmr_registers(1)(275) and tmr_registers(2)(275)) or                                                       
                            (tmr_registers(0)(275) and tmr_registers(2)(275));                                                         
                                                                                                                                     
        global_tmr_voter(0)(276)  <=    (tmr_registers(0)(276) and tmr_registers(1)(276)) or                                            
                            (tmr_registers(1)(276) and tmr_registers(2)(276)) or                                                       
                            (tmr_registers(0)(276) and tmr_registers(2)(276));                                                         
                                                                                                                                     
        global_tmr_voter(0)(277)  <=    (tmr_registers(0)(277) and tmr_registers(1)(277)) or                                            
                            (tmr_registers(1)(277) and tmr_registers(2)(277)) or                                                       
                            (tmr_registers(0)(277) and tmr_registers(2)(277));                                                         
                                                                                                                                     
        global_tmr_voter(0)(278)  <=    (tmr_registers(0)(278) and tmr_registers(1)(278)) or                                            
                            (tmr_registers(1)(278) and tmr_registers(2)(278)) or                                                       
                            (tmr_registers(0)(278) and tmr_registers(2)(278));                                                         
                                                                                                                                     
        global_tmr_voter(0)(279)  <=    (tmr_registers(0)(279) and tmr_registers(1)(279)) or                                            
                            (tmr_registers(1)(279) and tmr_registers(2)(279)) or                                                       
                            (tmr_registers(0)(279) and tmr_registers(2)(279));                                                         
                                                                                                                                     
        global_tmr_voter(0)(280)  <=    (tmr_registers(0)(280) and tmr_registers(1)(280)) or                                            
                            (tmr_registers(1)(280) and tmr_registers(2)(280)) or                                                       
                            (tmr_registers(0)(280) and tmr_registers(2)(280));                                                         
                                                                                                                                     
        global_tmr_voter(0)(281)  <=    (tmr_registers(0)(281) and tmr_registers(1)(281)) or                                            
                            (tmr_registers(1)(281) and tmr_registers(2)(281)) or                                                       
                            (tmr_registers(0)(281) and tmr_registers(2)(281));                                                         
                                                                                                                                     
        global_tmr_voter(0)(282)  <=    (tmr_registers(0)(282) and tmr_registers(1)(282)) or                                            
                            (tmr_registers(1)(282) and tmr_registers(2)(282)) or                                                       
                            (tmr_registers(0)(282) and tmr_registers(2)(282));                                                         
                                                                                                                                     
        global_tmr_voter(0)(283)  <=    (tmr_registers(0)(283) and tmr_registers(1)(283)) or                                            
                            (tmr_registers(1)(283) and tmr_registers(2)(283)) or                                                       
                            (tmr_registers(0)(283) and tmr_registers(2)(283));                                                         
                                                                                                                                     
        global_tmr_voter(0)(284)  <=    (tmr_registers(0)(284) and tmr_registers(1)(284)) or                                            
                            (tmr_registers(1)(284) and tmr_registers(2)(284)) or                                                       
                            (tmr_registers(0)(284) and tmr_registers(2)(284));                                                         
                                                                                                                                     
        global_tmr_voter(0)(285)  <=    (tmr_registers(0)(285) and tmr_registers(1)(285)) or                                            
                            (tmr_registers(1)(285) and tmr_registers(2)(285)) or                                                       
                            (tmr_registers(0)(285) and tmr_registers(2)(285));                                                         
                                                                                                                                     
        global_tmr_voter(0)(286)  <=    (tmr_registers(0)(286) and tmr_registers(1)(286)) or                                            
                            (tmr_registers(1)(286) and tmr_registers(2)(286)) or                                                       
                            (tmr_registers(0)(286) and tmr_registers(2)(286));                                                         
                                                                                                                                     
        global_tmr_voter(0)(287)  <=    (tmr_registers(0)(287) and tmr_registers(1)(287)) or                                            
                            (tmr_registers(1)(287) and tmr_registers(2)(287)) or                                                       
                            (tmr_registers(0)(287) and tmr_registers(2)(287));                                                         
                                                                                                                                     
        global_tmr_voter(0)(288)  <=    (tmr_registers(0)(288) and tmr_registers(1)(288)) or                                            
                            (tmr_registers(1)(288) and tmr_registers(2)(288)) or                                                       
                            (tmr_registers(0)(288) and tmr_registers(2)(288));                                                         
                                                                                                                                     
        global_tmr_voter(0)(289)  <=    (tmr_registers(0)(289) and tmr_registers(1)(289)) or                                            
                            (tmr_registers(1)(289) and tmr_registers(2)(289)) or                                                       
                            (tmr_registers(0)(289) and tmr_registers(2)(289));                                                         
                                                                                                                                     
        global_tmr_voter(0)(290)  <=    (tmr_registers(0)(290) and tmr_registers(1)(290)) or                                            
                            (tmr_registers(1)(290) and tmr_registers(2)(290)) or                                                       
                            (tmr_registers(0)(290) and tmr_registers(2)(290));                                                         
                                                                                                                                     
        global_tmr_voter(0)(291)  <=    (tmr_registers(0)(291) and tmr_registers(1)(291)) or                                            
                            (tmr_registers(1)(291) and tmr_registers(2)(291)) or                                                       
                            (tmr_registers(0)(291) and tmr_registers(2)(291));                                                         
                                                                                                                                     
        global_tmr_voter(0)(292)  <=    (tmr_registers(0)(292) and tmr_registers(1)(292)) or                                            
                            (tmr_registers(1)(292) and tmr_registers(2)(292)) or                                                       
                            (tmr_registers(0)(292) and tmr_registers(2)(292));                                                         
                                                                                                                                     
        global_tmr_voter(0)(293)  <=    (tmr_registers(0)(293) and tmr_registers(1)(293)) or                                            
                            (tmr_registers(1)(293) and tmr_registers(2)(293)) or                                                       
                            (tmr_registers(0)(293) and tmr_registers(2)(293));                                                         
                                                                                                                                     
        global_tmr_voter(0)(294)  <=    (tmr_registers(0)(294) and tmr_registers(1)(294)) or                                            
                            (tmr_registers(1)(294) and tmr_registers(2)(294)) or                                                       
                            (tmr_registers(0)(294) and tmr_registers(2)(294));                                                         
                                                                                                                                     
        global_tmr_voter(0)(295)  <=    (tmr_registers(0)(295) and tmr_registers(1)(295)) or                                            
                            (tmr_registers(1)(295) and tmr_registers(2)(295)) or                                                       
                            (tmr_registers(0)(295) and tmr_registers(2)(295));                                                         
                                                                                                                                     
        global_tmr_voter(0)(296)  <=    (tmr_registers(0)(296) and tmr_registers(1)(296)) or                                            
                            (tmr_registers(1)(296) and tmr_registers(2)(296)) or                                                       
                            (tmr_registers(0)(296) and tmr_registers(2)(296));                                                         
                                                                                                                                     
        global_tmr_voter(0)(297)  <=    (tmr_registers(0)(297) and tmr_registers(1)(297)) or                                            
                            (tmr_registers(1)(297) and tmr_registers(2)(297)) or                                                       
                            (tmr_registers(0)(297) and tmr_registers(2)(297));                                                         
                                                                                                                                     
        global_tmr_voter(0)(298)  <=    (tmr_registers(0)(298) and tmr_registers(1)(298)) or                                            
                            (tmr_registers(1)(298) and tmr_registers(2)(298)) or                                                       
                            (tmr_registers(0)(298) and tmr_registers(2)(298));                                                         
                                                                                                                                     
        global_tmr_voter(0)(299)  <=    (tmr_registers(0)(299) and tmr_registers(1)(299)) or                                            
                            (tmr_registers(1)(299) and tmr_registers(2)(299)) or                                                       
                            (tmr_registers(0)(299) and tmr_registers(2)(299));                                                         
                                                                                                                                     
        global_tmr_voter(0)(300)  <=    (tmr_registers(0)(300) and tmr_registers(1)(300)) or                                            
                            (tmr_registers(1)(300) and tmr_registers(2)(300)) or                                                       
                            (tmr_registers(0)(300) and tmr_registers(2)(300));                                                         
                                                                                                                                     
        global_tmr_voter(0)(301)  <=    (tmr_registers(0)(301) and tmr_registers(1)(301)) or                                            
                            (tmr_registers(1)(301) and tmr_registers(2)(301)) or                                                       
                            (tmr_registers(0)(301) and tmr_registers(2)(301));                                                         
                                                                                                                                     
        global_tmr_voter(0)(302)  <=    (tmr_registers(0)(302) and tmr_registers(1)(302)) or                                            
                            (tmr_registers(1)(302) and tmr_registers(2)(302)) or                                                       
                            (tmr_registers(0)(302) and tmr_registers(2)(302));                                                         
                                                                                                                                     
        global_tmr_voter(0)(303)  <=    (tmr_registers(0)(303) and tmr_registers(1)(303)) or                                            
                            (tmr_registers(1)(303) and tmr_registers(2)(303)) or                                                       
                            (tmr_registers(0)(303) and tmr_registers(2)(303));                                                         
                                                                                                                                     
        global_tmr_voter(0)(304)  <=    (tmr_registers(0)(304) and tmr_registers(1)(304)) or                                            
                            (tmr_registers(1)(304) and tmr_registers(2)(304)) or                                                       
                            (tmr_registers(0)(304) and tmr_registers(2)(304));                                                         
                                                                                                                                     
        global_tmr_voter(0)(305)  <=    (tmr_registers(0)(305) and tmr_registers(1)(305)) or                                            
                            (tmr_registers(1)(305) and tmr_registers(2)(305)) or                                                       
                            (tmr_registers(0)(305) and tmr_registers(2)(305));                                                         
                                                                                                                                     
        global_tmr_voter(0)(306)  <=    (tmr_registers(0)(306) and tmr_registers(1)(306)) or                                            
                            (tmr_registers(1)(306) and tmr_registers(2)(306)) or                                                       
                            (tmr_registers(0)(306) and tmr_registers(2)(306));                                                         
                                                                                                                                     
        global_tmr_voter(0)(307)  <=    (tmr_registers(0)(307) and tmr_registers(1)(307)) or                                            
                            (tmr_registers(1)(307) and tmr_registers(2)(307)) or                                                       
                            (tmr_registers(0)(307) and tmr_registers(2)(307));                                                         
                                                                                                                                     
        global_tmr_voter(0)(308)  <=    (tmr_registers(0)(308) and tmr_registers(1)(308)) or                                            
                            (tmr_registers(1)(308) and tmr_registers(2)(308)) or                                                       
                            (tmr_registers(0)(308) and tmr_registers(2)(308));                                                         
                                                                                                                                     
        global_tmr_voter(0)(309)  <=    (tmr_registers(0)(309) and tmr_registers(1)(309)) or                                            
                            (tmr_registers(1)(309) and tmr_registers(2)(309)) or                                                       
                            (tmr_registers(0)(309) and tmr_registers(2)(309));                                                         
                                                                                                                                     
        global_tmr_voter(0)(310)  <=    (tmr_registers(0)(310) and tmr_registers(1)(310)) or                                            
                            (tmr_registers(1)(310) and tmr_registers(2)(310)) or                                                       
                            (tmr_registers(0)(310) and tmr_registers(2)(310));                                                         
                                                                                                                                     
        global_tmr_voter(0)(311)  <=    (tmr_registers(0)(311) and tmr_registers(1)(311)) or                                            
                            (tmr_registers(1)(311) and tmr_registers(2)(311)) or                                                       
                            (tmr_registers(0)(311) and tmr_registers(2)(311));                                                         
                                                                                                                                     
        global_tmr_voter(0)(312)  <=    (tmr_registers(0)(312) and tmr_registers(1)(312)) or                                            
                            (tmr_registers(1)(312) and tmr_registers(2)(312)) or                                                       
                            (tmr_registers(0)(312) and tmr_registers(2)(312));                                                         
                                                                                                                                     
        global_tmr_voter(0)(313)  <=    (tmr_registers(0)(313) and tmr_registers(1)(313)) or                                            
                            (tmr_registers(1)(313) and tmr_registers(2)(313)) or                                                       
                            (tmr_registers(0)(313) and tmr_registers(2)(313));                                                         
                                                                                                                                     
        global_tmr_voter(0)(314)  <=    (tmr_registers(0)(314) and tmr_registers(1)(314)) or                                            
                            (tmr_registers(1)(314) and tmr_registers(2)(314)) or                                                       
                            (tmr_registers(0)(314) and tmr_registers(2)(314));                                                         
                                                                                                                                     
        global_tmr_voter(0)(315)  <=    (tmr_registers(0)(315) and tmr_registers(1)(315)) or                                            
                            (tmr_registers(1)(315) and tmr_registers(2)(315)) or                                                       
                            (tmr_registers(0)(315) and tmr_registers(2)(315));                                                         
                                                                                                                                     
        global_tmr_voter(0)(316)  <=    (tmr_registers(0)(316) and tmr_registers(1)(316)) or                                            
                            (tmr_registers(1)(316) and tmr_registers(2)(316)) or                                                       
                            (tmr_registers(0)(316) and tmr_registers(2)(316));                                                         
                                                                                                                                     
        global_tmr_voter(0)(317)  <=    (tmr_registers(0)(317) and tmr_registers(1)(317)) or                                            
                            (tmr_registers(1)(317) and tmr_registers(2)(317)) or                                                       
                            (tmr_registers(0)(317) and tmr_registers(2)(317));                                                         
                                                                                                                                     
        global_tmr_voter(0)(318)  <=    (tmr_registers(0)(318) and tmr_registers(1)(318)) or                                            
                            (tmr_registers(1)(318) and tmr_registers(2)(318)) or                                                       
                            (tmr_registers(0)(318) and tmr_registers(2)(318));                                                         
                                                                                                                                     
        global_tmr_voter(0)(319)  <=    (tmr_registers(0)(319) and tmr_registers(1)(319)) or                                            
                            (tmr_registers(1)(319) and tmr_registers(2)(319)) or                                                       
                            (tmr_registers(0)(319) and tmr_registers(2)(319));                                                         
                                                                                                                                     
        global_tmr_voter(0)(320)  <=    (tmr_registers(0)(320) and tmr_registers(1)(320)) or                                            
                            (tmr_registers(1)(320) and tmr_registers(2)(320)) or                                                       
                            (tmr_registers(0)(320) and tmr_registers(2)(320));                                                         
                                                                                                                                     
        global_tmr_voter(0)(321)  <=    (tmr_registers(0)(321) and tmr_registers(1)(321)) or                                            
                            (tmr_registers(1)(321) and tmr_registers(2)(321)) or                                                       
                            (tmr_registers(0)(321) and tmr_registers(2)(321));                                                         
                                                                                                                                     
        global_tmr_voter(0)(322)  <=    (tmr_registers(0)(322) and tmr_registers(1)(322)) or                                            
                            (tmr_registers(1)(322) and tmr_registers(2)(322)) or                                                       
                            (tmr_registers(0)(322) and tmr_registers(2)(322));                                                         
                                                                                                                                     
        global_tmr_voter(0)(323)  <=    (tmr_registers(0)(323) and tmr_registers(1)(323)) or                                            
                            (tmr_registers(1)(323) and tmr_registers(2)(323)) or                                                       
                            (tmr_registers(0)(323) and tmr_registers(2)(323));                                                         
                                                                                                                                     
        global_tmr_voter(0)(324)  <=    (tmr_registers(0)(324) and tmr_registers(1)(324)) or                                            
                            (tmr_registers(1)(324) and tmr_registers(2)(324)) or                                                       
                            (tmr_registers(0)(324) and tmr_registers(2)(324));                                                         
                                                                                                                                     
        global_tmr_voter(0)(325)  <=    (tmr_registers(0)(325) and tmr_registers(1)(325)) or                                            
                            (tmr_registers(1)(325) and tmr_registers(2)(325)) or                                                       
                            (tmr_registers(0)(325) and tmr_registers(2)(325));                                                         
                                                                                                                                     
        global_tmr_voter(0)(326)  <=    (tmr_registers(0)(326) and tmr_registers(1)(326)) or                                            
                            (tmr_registers(1)(326) and tmr_registers(2)(326)) or                                                       
                            (tmr_registers(0)(326) and tmr_registers(2)(326));                                                         
                                                                                                                                     
        global_tmr_voter(0)(327)  <=    (tmr_registers(0)(327) and tmr_registers(1)(327)) or                                            
                            (tmr_registers(1)(327) and tmr_registers(2)(327)) or                                                       
                            (tmr_registers(0)(327) and tmr_registers(2)(327));                                                         
                                                                                                                                     
        global_tmr_voter(0)(328)  <=    (tmr_registers(0)(328) and tmr_registers(1)(328)) or                                            
                            (tmr_registers(1)(328) and tmr_registers(2)(328)) or                                                       
                            (tmr_registers(0)(328) and tmr_registers(2)(328));                                                         
                                                                                                                                     
        global_tmr_voter(0)(329)  <=    (tmr_registers(0)(329) and tmr_registers(1)(329)) or                                            
                            (tmr_registers(1)(329) and tmr_registers(2)(329)) or                                                       
                            (tmr_registers(0)(329) and tmr_registers(2)(329));                                                         
                                                                                                                                     
        global_tmr_voter(0)(330)  <=    (tmr_registers(0)(330) and tmr_registers(1)(330)) or                                            
                            (tmr_registers(1)(330) and tmr_registers(2)(330)) or                                                       
                            (tmr_registers(0)(330) and tmr_registers(2)(330));                                                         
                                                                                                                                     
        global_tmr_voter(0)(331)  <=    (tmr_registers(0)(331) and tmr_registers(1)(331)) or                                            
                            (tmr_registers(1)(331) and tmr_registers(2)(331)) or                                                       
                            (tmr_registers(0)(331) and tmr_registers(2)(331));                                                         
                                                                                                                                     
        global_tmr_voter(0)(332)  <=    (tmr_registers(0)(332) and tmr_registers(1)(332)) or                                            
                            (tmr_registers(1)(332) and tmr_registers(2)(332)) or                                                       
                            (tmr_registers(0)(332) and tmr_registers(2)(332));                                                         
                                                                                                                                     
        global_tmr_voter(0)(333)  <=    (tmr_registers(0)(333) and tmr_registers(1)(333)) or                                            
                            (tmr_registers(1)(333) and tmr_registers(2)(333)) or                                                       
                            (tmr_registers(0)(333) and tmr_registers(2)(333));                                                         
                                                                                                                                     
        global_tmr_voter(0)(334)  <=    (tmr_registers(0)(334) and tmr_registers(1)(334)) or                                            
                            (tmr_registers(1)(334) and tmr_registers(2)(334)) or                                                       
                            (tmr_registers(0)(334) and tmr_registers(2)(334));                                                         
                                                                                                                                     
        global_tmr_voter(0)(335)  <=    (tmr_registers(0)(335) and tmr_registers(1)(335)) or                                            
                            (tmr_registers(1)(335) and tmr_registers(2)(335)) or                                                       
                            (tmr_registers(0)(335) and tmr_registers(2)(335));                                                         
                                                                                                                                     
        global_tmr_voter(0)(336)  <=    (tmr_registers(0)(336) and tmr_registers(1)(336)) or                                            
                            (tmr_registers(1)(336) and tmr_registers(2)(336)) or                                                       
                            (tmr_registers(0)(336) and tmr_registers(2)(336));                                                         
                                                                                                                                     
        global_tmr_voter(0)(337)  <=    (tmr_registers(0)(337) and tmr_registers(1)(337)) or                                            
                            (tmr_registers(1)(337) and tmr_registers(2)(337)) or                                                       
                            (tmr_registers(0)(337) and tmr_registers(2)(337));                                                         
                                                                                                                                     
        global_tmr_voter(0)(338)  <=    (tmr_registers(0)(338) and tmr_registers(1)(338)) or                                            
                            (tmr_registers(1)(338) and tmr_registers(2)(338)) or                                                       
                            (tmr_registers(0)(338) and tmr_registers(2)(338));                                                         
                                                                                                                                     
        global_tmr_voter(0)(339)  <=    (tmr_registers(0)(339) and tmr_registers(1)(339)) or                                            
                            (tmr_registers(1)(339) and tmr_registers(2)(339)) or                                                       
                            (tmr_registers(0)(339) and tmr_registers(2)(339));                                                         
                                                                                                                                     
        global_tmr_voter(0)(340)  <=    (tmr_registers(0)(340) and tmr_registers(1)(340)) or                                            
                            (tmr_registers(1)(340) and tmr_registers(2)(340)) or                                                       
                            (tmr_registers(0)(340) and tmr_registers(2)(340));                                                         
                                                                                                                                     
        global_tmr_voter(0)(341)  <=    (tmr_registers(0)(341) and tmr_registers(1)(341)) or                                            
                            (tmr_registers(1)(341) and tmr_registers(2)(341)) or                                                       
                            (tmr_registers(0)(341) and tmr_registers(2)(341));                                                         
                                                                                                                                     
        global_tmr_voter(0)(342)  <=    (tmr_registers(0)(342) and tmr_registers(1)(342)) or                                            
                            (tmr_registers(1)(342) and tmr_registers(2)(342)) or                                                       
                            (tmr_registers(0)(342) and tmr_registers(2)(342));                                                         
                                                                                                                                     
        global_tmr_voter(0)(343)  <=    (tmr_registers(0)(343) and tmr_registers(1)(343)) or                                            
                            (tmr_registers(1)(343) and tmr_registers(2)(343)) or                                                       
                            (tmr_registers(0)(343) and tmr_registers(2)(343));                                                         
                                                                                                                                     
        global_tmr_voter(0)(344)  <=    (tmr_registers(0)(344) and tmr_registers(1)(344)) or                                            
                            (tmr_registers(1)(344) and tmr_registers(2)(344)) or                                                       
                            (tmr_registers(0)(344) and tmr_registers(2)(344));                                                         
                                                                                                                                     
        global_tmr_voter(0)(345)  <=    (tmr_registers(0)(345) and tmr_registers(1)(345)) or                                            
                            (tmr_registers(1)(345) and tmr_registers(2)(345)) or                                                       
                            (tmr_registers(0)(345) and tmr_registers(2)(345));                                                         
                                                                                                                                     
        global_tmr_voter(0)(346)  <=    (tmr_registers(0)(346) and tmr_registers(1)(346)) or                                            
                            (tmr_registers(1)(346) and tmr_registers(2)(346)) or                                                       
                            (tmr_registers(0)(346) and tmr_registers(2)(346));                                                         
                                                                                                                                     
        global_tmr_voter(0)(347)  <=    (tmr_registers(0)(347) and tmr_registers(1)(347)) or                                            
                            (tmr_registers(1)(347) and tmr_registers(2)(347)) or                                                       
                            (tmr_registers(0)(347) and tmr_registers(2)(347));                                                         
                                                                                                                                     
        global_tmr_voter(0)(348)  <=    (tmr_registers(0)(348) and tmr_registers(1)(348)) or                                            
                            (tmr_registers(1)(348) and tmr_registers(2)(348)) or                                                       
                            (tmr_registers(0)(348) and tmr_registers(2)(348));                                                         
                                                                                                                                     
        global_tmr_voter(0)(349)  <=    (tmr_registers(0)(349) and tmr_registers(1)(349)) or                                            
                            (tmr_registers(1)(349) and tmr_registers(2)(349)) or                                                       
                            (tmr_registers(0)(349) and tmr_registers(2)(349));                                                         
                                                                                                                                     
        global_tmr_voter(0)(350)  <=    (tmr_registers(0)(350) and tmr_registers(1)(350)) or                                            
                            (tmr_registers(1)(350) and tmr_registers(2)(350)) or                                                       
                            (tmr_registers(0)(350) and tmr_registers(2)(350));                                                         
                                                                                                                                     
        global_tmr_voter(0)(351)  <=    (tmr_registers(0)(351) and tmr_registers(1)(351)) or                                            
                            (tmr_registers(1)(351) and tmr_registers(2)(351)) or                                                       
                            (tmr_registers(0)(351) and tmr_registers(2)(351));                                                         
                                                                                                                                     
        global_tmr_voter(0)(352)  <=    (tmr_registers(0)(352) and tmr_registers(1)(352)) or                                            
                            (tmr_registers(1)(352) and tmr_registers(2)(352)) or                                                       
                            (tmr_registers(0)(352) and tmr_registers(2)(352));                                                         
                                                                                                                                     
        global_tmr_voter(0)(353)  <=    (tmr_registers(0)(353) and tmr_registers(1)(353)) or                                            
                            (tmr_registers(1)(353) and tmr_registers(2)(353)) or                                                       
                            (tmr_registers(0)(353) and tmr_registers(2)(353));                                                         
                                                                                                                                     
        global_tmr_voter(0)(354)  <=    (tmr_registers(0)(354) and tmr_registers(1)(354)) or                                            
                            (tmr_registers(1)(354) and tmr_registers(2)(354)) or                                                       
                            (tmr_registers(0)(354) and tmr_registers(2)(354));                                                         
                                                                                                                                     
        global_tmr_voter(0)(355)  <=    (tmr_registers(0)(355) and tmr_registers(1)(355)) or                                            
                            (tmr_registers(1)(355) and tmr_registers(2)(355)) or                                                       
                            (tmr_registers(0)(355) and tmr_registers(2)(355));                                                         
                                                                                                                                     
        global_tmr_voter(0)(356)  <=    (tmr_registers(0)(356) and tmr_registers(1)(356)) or                                            
                            (tmr_registers(1)(356) and tmr_registers(2)(356)) or                                                       
                            (tmr_registers(0)(356) and tmr_registers(2)(356));                                                         
                                                                                                                                     
        global_tmr_voter(0)(357)  <=    (tmr_registers(0)(357) and tmr_registers(1)(357)) or                                            
                            (tmr_registers(1)(357) and tmr_registers(2)(357)) or                                                       
                            (tmr_registers(0)(357) and tmr_registers(2)(357));                                                         
                                                                                                                                     
        global_tmr_voter(0)(358)  <=    (tmr_registers(0)(358) and tmr_registers(1)(358)) or                                            
                            (tmr_registers(1)(358) and tmr_registers(2)(358)) or                                                       
                            (tmr_registers(0)(358) and tmr_registers(2)(358));                                                         
                                                                                                                                     
        global_tmr_voter(0)(359)  <=    (tmr_registers(0)(359) and tmr_registers(1)(359)) or                                            
                            (tmr_registers(1)(359) and tmr_registers(2)(359)) or                                                       
                            (tmr_registers(0)(359) and tmr_registers(2)(359));                                                         
                                                                                                                                     
        global_tmr_voter(0)(360)  <=    (tmr_registers(0)(360) and tmr_registers(1)(360)) or                                            
                            (tmr_registers(1)(360) and tmr_registers(2)(360)) or                                                       
                            (tmr_registers(0)(360) and tmr_registers(2)(360));                                                         
                                                                                                                                     
        global_tmr_voter(0)(361)  <=    (tmr_registers(0)(361) and tmr_registers(1)(361)) or                                            
                            (tmr_registers(1)(361) and tmr_registers(2)(361)) or                                                       
                            (tmr_registers(0)(361) and tmr_registers(2)(361));                                                         
                                                                                                                                     
        global_tmr_voter(0)(362)  <=    (tmr_registers(0)(362) and tmr_registers(1)(362)) or                                            
                            (tmr_registers(1)(362) and tmr_registers(2)(362)) or                                                       
                            (tmr_registers(0)(362) and tmr_registers(2)(362));                                                         
                                                                                                                                     
        global_tmr_voter(0)(363)  <=    (tmr_registers(0)(363) and tmr_registers(1)(363)) or                                            
                            (tmr_registers(1)(363) and tmr_registers(2)(363)) or                                                       
                            (tmr_registers(0)(363) and tmr_registers(2)(363));                                                         
                                                                                                                                     
        global_tmr_voter(0)(364)  <=    (tmr_registers(0)(364) and tmr_registers(1)(364)) or                                            
                            (tmr_registers(1)(364) and tmr_registers(2)(364)) or                                                       
                            (tmr_registers(0)(364) and tmr_registers(2)(364));                                                         
                                                                                                                                     
        global_tmr_voter(0)(365)  <=    (tmr_registers(0)(365) and tmr_registers(1)(365)) or                                            
                            (tmr_registers(1)(365) and tmr_registers(2)(365)) or                                                       
                            (tmr_registers(0)(365) and tmr_registers(2)(365));                                                         
                                                                                                                                     
        global_tmr_voter(0)(366)  <=    (tmr_registers(0)(366) and tmr_registers(1)(366)) or                                            
                            (tmr_registers(1)(366) and tmr_registers(2)(366)) or                                                       
                            (tmr_registers(0)(366) and tmr_registers(2)(366));                                                         
                                                                                                                                     
        global_tmr_voter(0)(367)  <=    (tmr_registers(0)(367) and tmr_registers(1)(367)) or                                            
                            (tmr_registers(1)(367) and tmr_registers(2)(367)) or                                                       
                            (tmr_registers(0)(367) and tmr_registers(2)(367));                                                         
                                                                                                                                     
        global_tmr_voter(0)(368)  <=    (tmr_registers(0)(368) and tmr_registers(1)(368)) or                                            
                            (tmr_registers(1)(368) and tmr_registers(2)(368)) or                                                       
                            (tmr_registers(0)(368) and tmr_registers(2)(368));                                                         
                                                                                                                                     
        global_tmr_voter(0)(369)  <=    (tmr_registers(0)(369) and tmr_registers(1)(369)) or                                            
                            (tmr_registers(1)(369) and tmr_registers(2)(369)) or                                                       
                            (tmr_registers(0)(369) and tmr_registers(2)(369));                                                         
                                                                                                                                     
        global_tmr_voter(0)(370)  <=    (tmr_registers(0)(370) and tmr_registers(1)(370)) or                                            
                            (tmr_registers(1)(370) and tmr_registers(2)(370)) or                                                       
                            (tmr_registers(0)(370) and tmr_registers(2)(370));                                                         
                                                                                                                                     
        global_tmr_voter(0)(371)  <=    (tmr_registers(0)(371) and tmr_registers(1)(371)) or                                            
                            (tmr_registers(1)(371) and tmr_registers(2)(371)) or                                                       
                            (tmr_registers(0)(371) and tmr_registers(2)(371));                                                         
                                                                                                                                     
        global_tmr_voter(0)(372)  <=    (tmr_registers(0)(372) and tmr_registers(1)(372)) or                                            
                            (tmr_registers(1)(372) and tmr_registers(2)(372)) or                                                       
                            (tmr_registers(0)(372) and tmr_registers(2)(372));                                                         
                                                                                                                                     
        global_tmr_voter(0)(373)  <=    (tmr_registers(0)(373) and tmr_registers(1)(373)) or                                            
                            (tmr_registers(1)(373) and tmr_registers(2)(373)) or                                                       
                            (tmr_registers(0)(373) and tmr_registers(2)(373));                                                         
                                                                                                                                     
        global_tmr_voter(0)(374)  <=    (tmr_registers(0)(374) and tmr_registers(1)(374)) or                                            
                            (tmr_registers(1)(374) and tmr_registers(2)(374)) or                                                       
                            (tmr_registers(0)(374) and tmr_registers(2)(374));                                                         
                                                                                                                                     
        global_tmr_voter(0)(375)  <=    (tmr_registers(0)(375) and tmr_registers(1)(375)) or                                            
                            (tmr_registers(1)(375) and tmr_registers(2)(375)) or                                                       
                            (tmr_registers(0)(375) and tmr_registers(2)(375));                                                         
                                                                                                                                     
        global_tmr_voter(0)(376)  <=    (tmr_registers(0)(376) and tmr_registers(1)(376)) or                                            
                            (tmr_registers(1)(376) and tmr_registers(2)(376)) or                                                       
                            (tmr_registers(0)(376) and tmr_registers(2)(376));                                                         
                                                                                                                                     
        global_tmr_voter(0)(377)  <=    (tmr_registers(0)(377) and tmr_registers(1)(377)) or                                            
                            (tmr_registers(1)(377) and tmr_registers(2)(377)) or                                                       
                            (tmr_registers(0)(377) and tmr_registers(2)(377));                                                         
                                                                                                                                     
        global_tmr_voter(0)(378)  <=    (tmr_registers(0)(378) and tmr_registers(1)(378)) or                                            
                            (tmr_registers(1)(378) and tmr_registers(2)(378)) or                                                       
                            (tmr_registers(0)(378) and tmr_registers(2)(378));                                                         
                                                                                                                                     
        global_tmr_voter(0)(379)  <=    (tmr_registers(0)(379) and tmr_registers(1)(379)) or                                            
                            (tmr_registers(1)(379) and tmr_registers(2)(379)) or                                                       
                            (tmr_registers(0)(379) and tmr_registers(2)(379));                                                         
                                                                                                                                     
        global_tmr_voter(0)(380)  <=    (tmr_registers(0)(380) and tmr_registers(1)(380)) or                                            
                            (tmr_registers(1)(380) and tmr_registers(2)(380)) or                                                       
                            (tmr_registers(0)(380) and tmr_registers(2)(380));                                                         
                                                                                                                                     
        global_tmr_voter(0)(381)  <=    (tmr_registers(0)(381) and tmr_registers(1)(381)) or                                            
                            (tmr_registers(1)(381) and tmr_registers(2)(381)) or                                                       
                            (tmr_registers(0)(381) and tmr_registers(2)(381));                                                         
                                                                                                                                     
        global_tmr_voter(0)(382)  <=    (tmr_registers(0)(382) and tmr_registers(1)(382)) or                                            
                            (tmr_registers(1)(382) and tmr_registers(2)(382)) or                                                       
                            (tmr_registers(0)(382) and tmr_registers(2)(382));                                                         
                                                                                                                                     
        global_tmr_voter(0)(383)  <=    (tmr_registers(0)(383) and tmr_registers(1)(383)) or                                            
                            (tmr_registers(1)(383) and tmr_registers(2)(383)) or                                                       
                            (tmr_registers(0)(383) and tmr_registers(2)(383));                                                         
                                                                                                                                     
        global_tmr_voter(0)(384)  <=    (tmr_registers(0)(384) and tmr_registers(1)(384)) or                                            
                            (tmr_registers(1)(384) and tmr_registers(2)(384)) or                                                       
                            (tmr_registers(0)(384) and tmr_registers(2)(384));                                                         
                                                                                                                                     
        global_tmr_voter(0)(385)  <=    (tmr_registers(0)(385) and tmr_registers(1)(385)) or                                            
                            (tmr_registers(1)(385) and tmr_registers(2)(385)) or                                                       
                            (tmr_registers(0)(385) and tmr_registers(2)(385));                                                         
                                                                                                                                     
        global_tmr_voter(0)(386)  <=    (tmr_registers(0)(386) and tmr_registers(1)(386)) or                                            
                            (tmr_registers(1)(386) and tmr_registers(2)(386)) or                                                       
                            (tmr_registers(0)(386) and tmr_registers(2)(386));                                                         
                                                                                                                                     
        global_tmr_voter(0)(387)  <=    (tmr_registers(0)(387) and tmr_registers(1)(387)) or                                            
                            (tmr_registers(1)(387) and tmr_registers(2)(387)) or                                                       
                            (tmr_registers(0)(387) and tmr_registers(2)(387));                                                         
                                                                                                                                     
        global_tmr_voter(0)(388)  <=    (tmr_registers(0)(388) and tmr_registers(1)(388)) or                                            
                            (tmr_registers(1)(388) and tmr_registers(2)(388)) or                                                       
                            (tmr_registers(0)(388) and tmr_registers(2)(388));                                                         
                                                                                                                                     
        global_tmr_voter(0)(389)  <=    (tmr_registers(0)(389) and tmr_registers(1)(389)) or                                            
                            (tmr_registers(1)(389) and tmr_registers(2)(389)) or                                                       
                            (tmr_registers(0)(389) and tmr_registers(2)(389));                                                         
                                                                                                                                     
        global_tmr_voter(0)(390)  <=    (tmr_registers(0)(390) and tmr_registers(1)(390)) or                                            
                            (tmr_registers(1)(390) and tmr_registers(2)(390)) or                                                       
                            (tmr_registers(0)(390) and tmr_registers(2)(390));                                                         
                                                                                                                                     
        global_tmr_voter(0)(391)  <=    (tmr_registers(0)(391) and tmr_registers(1)(391)) or                                            
                            (tmr_registers(1)(391) and tmr_registers(2)(391)) or                                                       
                            (tmr_registers(0)(391) and tmr_registers(2)(391));                                                         
                                                                                                                                     
        global_tmr_voter(0)(392)  <=    (tmr_registers(0)(392) and tmr_registers(1)(392)) or                                            
                            (tmr_registers(1)(392) and tmr_registers(2)(392)) or                                                       
                            (tmr_registers(0)(392) and tmr_registers(2)(392));                                                         
                                                                                                                                     
        global_tmr_voter(0)(393)  <=    (tmr_registers(0)(393) and tmr_registers(1)(393)) or                                            
                            (tmr_registers(1)(393) and tmr_registers(2)(393)) or                                                       
                            (tmr_registers(0)(393) and tmr_registers(2)(393));                                                         
                                                                                                                                     
        global_tmr_voter(0)(394)  <=    (tmr_registers(0)(394) and tmr_registers(1)(394)) or                                            
                            (tmr_registers(1)(394) and tmr_registers(2)(394)) or                                                       
                            (tmr_registers(0)(394) and tmr_registers(2)(394));                                                         
                                                                                                                                     
        global_tmr_voter(0)(395)  <=    (tmr_registers(0)(395) and tmr_registers(1)(395)) or                                            
                            (tmr_registers(1)(395) and tmr_registers(2)(395)) or                                                       
                            (tmr_registers(0)(395) and tmr_registers(2)(395));                                                         
                                                                                                                                     
        global_tmr_voter(0)(396)  <=    (tmr_registers(0)(396) and tmr_registers(1)(396)) or                                            
                            (tmr_registers(1)(396) and tmr_registers(2)(396)) or                                                       
                            (tmr_registers(0)(396) and tmr_registers(2)(396));                                                         
                                                                                                                                     
        global_tmr_voter(0)(397)  <=    (tmr_registers(0)(397) and tmr_registers(1)(397)) or                                            
                            (tmr_registers(1)(397) and tmr_registers(2)(397)) or                                                       
                            (tmr_registers(0)(397) and tmr_registers(2)(397));                                                         
                                                                                                                                     
        global_tmr_voter(0)(398)  <=    (tmr_registers(0)(398) and tmr_registers(1)(398)) or                                            
                            (tmr_registers(1)(398) and tmr_registers(2)(398)) or                                                       
                            (tmr_registers(0)(398) and tmr_registers(2)(398));                                                         
                                                                                                                                     
        global_tmr_voter(0)(399)  <=    (tmr_registers(0)(399) and tmr_registers(1)(399)) or                                            
                            (tmr_registers(1)(399) and tmr_registers(2)(399)) or                                                       
                            (tmr_registers(0)(399) and tmr_registers(2)(399));                                                         
                                                                                                                                     
        global_tmr_voter(0)(400)  <=    (tmr_registers(0)(400) and tmr_registers(1)(400)) or                                            
                            (tmr_registers(1)(400) and tmr_registers(2)(400)) or                                                       
                            (tmr_registers(0)(400) and tmr_registers(2)(400));                                                         
                                                                                                                                     
        global_tmr_voter(0)(401)  <=    (tmr_registers(0)(401) and tmr_registers(1)(401)) or                                            
                            (tmr_registers(1)(401) and tmr_registers(2)(401)) or                                                       
                            (tmr_registers(0)(401) and tmr_registers(2)(401));                                                         
                                                                                                                                     
        global_tmr_voter(0)(402)  <=    (tmr_registers(0)(402) and tmr_registers(1)(402)) or                                            
                            (tmr_registers(1)(402) and tmr_registers(2)(402)) or                                                       
                            (tmr_registers(0)(402) and tmr_registers(2)(402));                                                         
                                                                                                                                     
        global_tmr_voter(0)(403)  <=    (tmr_registers(0)(403) and tmr_registers(1)(403)) or                                            
                            (tmr_registers(1)(403) and tmr_registers(2)(403)) or                                                       
                            (tmr_registers(0)(403) and tmr_registers(2)(403));                                                         
                                                                                                                                     
        global_tmr_voter(0)(404)  <=    (tmr_registers(0)(404) and tmr_registers(1)(404)) or                                            
                            (tmr_registers(1)(404) and tmr_registers(2)(404)) or                                                       
                            (tmr_registers(0)(404) and tmr_registers(2)(404));                                                         
                                                                                                                                     
        global_tmr_voter(0)(405)  <=    (tmr_registers(0)(405) and tmr_registers(1)(405)) or                                            
                            (tmr_registers(1)(405) and tmr_registers(2)(405)) or                                                       
                            (tmr_registers(0)(405) and tmr_registers(2)(405));                                                         
                                                                                                                                     
        global_tmr_voter(0)(406)  <=    (tmr_registers(0)(406) and tmr_registers(1)(406)) or                                            
                            (tmr_registers(1)(406) and tmr_registers(2)(406)) or                                                       
                            (tmr_registers(0)(406) and tmr_registers(2)(406));                                                         
                                                                                                                                     
        global_tmr_voter(0)(407)  <=    (tmr_registers(0)(407) and tmr_registers(1)(407)) or                                            
                            (tmr_registers(1)(407) and tmr_registers(2)(407)) or                                                       
                            (tmr_registers(0)(407) and tmr_registers(2)(407));                                                         
                                                                                                                                     
        global_tmr_voter(0)(408)  <=    (tmr_registers(0)(408) and tmr_registers(1)(408)) or                                            
                            (tmr_registers(1)(408) and tmr_registers(2)(408)) or                                                       
                            (tmr_registers(0)(408) and tmr_registers(2)(408));                                                         
                                                                                                                                     
        global_tmr_voter(0)(409)  <=    (tmr_registers(0)(409) and tmr_registers(1)(409)) or                                            
                            (tmr_registers(1)(409) and tmr_registers(2)(409)) or                                                       
                            (tmr_registers(0)(409) and tmr_registers(2)(409));                                                         
                                                                                                                                     
        global_tmr_voter(0)(410)  <=    (tmr_registers(0)(410) and tmr_registers(1)(410)) or                                            
                            (tmr_registers(1)(410) and tmr_registers(2)(410)) or                                                       
                            (tmr_registers(0)(410) and tmr_registers(2)(410));                                                         
                                                                                                                                     
        global_tmr_voter(0)(411)  <=    (tmr_registers(0)(411) and tmr_registers(1)(411)) or                                            
                            (tmr_registers(1)(411) and tmr_registers(2)(411)) or                                                       
                            (tmr_registers(0)(411) and tmr_registers(2)(411));                                                         
                                                                                                                                     
        global_tmr_voter(0)(412)  <=    (tmr_registers(0)(412) and tmr_registers(1)(412)) or                                            
                            (tmr_registers(1)(412) and tmr_registers(2)(412)) or                                                       
                            (tmr_registers(0)(412) and tmr_registers(2)(412));                                                         
                                                                                                                                     
        global_tmr_voter(0)(413)  <=    (tmr_registers(0)(413) and tmr_registers(1)(413)) or                                            
                            (tmr_registers(1)(413) and tmr_registers(2)(413)) or                                                       
                            (tmr_registers(0)(413) and tmr_registers(2)(413));                                                         
                                                                                                                                     
        global_tmr_voter(0)(414)  <=    (tmr_registers(0)(414) and tmr_registers(1)(414)) or                                            
                            (tmr_registers(1)(414) and tmr_registers(2)(414)) or                                                       
                            (tmr_registers(0)(414) and tmr_registers(2)(414));                                                         
                                                                                                                                     
        global_tmr_voter(0)(415)  <=    (tmr_registers(0)(415) and tmr_registers(1)(415)) or                                            
                            (tmr_registers(1)(415) and tmr_registers(2)(415)) or                                                       
                            (tmr_registers(0)(415) and tmr_registers(2)(415));                                                         
                                                                                                                                     
        global_tmr_voter(0)(416)  <=    (tmr_registers(0)(416) and tmr_registers(1)(416)) or                                            
                            (tmr_registers(1)(416) and tmr_registers(2)(416)) or                                                       
                            (tmr_registers(0)(416) and tmr_registers(2)(416));                                                         
                                                                                                                                     
        global_tmr_voter(0)(417)  <=    (tmr_registers(0)(417) and tmr_registers(1)(417)) or                                            
                            (tmr_registers(1)(417) and tmr_registers(2)(417)) or                                                       
                            (tmr_registers(0)(417) and tmr_registers(2)(417));                                                         
                                                                                                                                     
        global_tmr_voter(0)(418)  <=    (tmr_registers(0)(418) and tmr_registers(1)(418)) or                                            
                            (tmr_registers(1)(418) and tmr_registers(2)(418)) or                                                       
                            (tmr_registers(0)(418) and tmr_registers(2)(418));                                                         
                                                                                                                                     
        global_tmr_voter(0)(419)  <=    (tmr_registers(0)(419) and tmr_registers(1)(419)) or                                            
                            (tmr_registers(1)(419) and tmr_registers(2)(419)) or                                                       
                            (tmr_registers(0)(419) and tmr_registers(2)(419));                                                         
                                                                                                                                     
        global_tmr_voter(0)(420)  <=    (tmr_registers(0)(420) and tmr_registers(1)(420)) or                                            
                            (tmr_registers(1)(420) and tmr_registers(2)(420)) or                                                       
                            (tmr_registers(0)(420) and tmr_registers(2)(420));                                                         
                                                                                                                                     
        global_tmr_voter(0)(421)  <=    (tmr_registers(0)(421) and tmr_registers(1)(421)) or                                            
                            (tmr_registers(1)(421) and tmr_registers(2)(421)) or                                                       
                            (tmr_registers(0)(421) and tmr_registers(2)(421));                                                         
                                                                                                                                     
        global_tmr_voter(0)(422)  <=    (tmr_registers(0)(422) and tmr_registers(1)(422)) or                                            
                            (tmr_registers(1)(422) and tmr_registers(2)(422)) or                                                       
                            (tmr_registers(0)(422) and tmr_registers(2)(422));                                                         
                                                                                                                                     
        global_tmr_voter(0)(423)  <=    (tmr_registers(0)(423) and tmr_registers(1)(423)) or                                            
                            (tmr_registers(1)(423) and tmr_registers(2)(423)) or                                                       
                            (tmr_registers(0)(423) and tmr_registers(2)(423));                                                         
                                                                                                                                     
        global_tmr_voter(0)(424)  <=    (tmr_registers(0)(424) and tmr_registers(1)(424)) or                                            
                            (tmr_registers(1)(424) and tmr_registers(2)(424)) or                                                       
                            (tmr_registers(0)(424) and tmr_registers(2)(424));                                                         
                                                                                                                                     
        global_tmr_voter(0)(425)  <=    (tmr_registers(0)(425) and tmr_registers(1)(425)) or                                            
                            (tmr_registers(1)(425) and tmr_registers(2)(425)) or                                                       
                            (tmr_registers(0)(425) and tmr_registers(2)(425));                                                         
                                                                                                                                     
        global_tmr_voter(0)(426)  <=    (tmr_registers(0)(426) and tmr_registers(1)(426)) or                                            
                            (tmr_registers(1)(426) and tmr_registers(2)(426)) or                                                       
                            (tmr_registers(0)(426) and tmr_registers(2)(426));                                                         
                                                                                                                                     
        global_tmr_voter(0)(427)  <=    (tmr_registers(0)(427) and tmr_registers(1)(427)) or                                            
                            (tmr_registers(1)(427) and tmr_registers(2)(427)) or                                                       
                            (tmr_registers(0)(427) and tmr_registers(2)(427));                                                         
                                                                                                                                     
        global_tmr_voter(0)(428)  <=    (tmr_registers(0)(428) and tmr_registers(1)(428)) or                                            
                            (tmr_registers(1)(428) and tmr_registers(2)(428)) or                                                       
                            (tmr_registers(0)(428) and tmr_registers(2)(428));                                                         
                                                                                                                                     
        global_tmr_voter(0)(429)  <=    (tmr_registers(0)(429) and tmr_registers(1)(429)) or                                            
                            (tmr_registers(1)(429) and tmr_registers(2)(429)) or                                                       
                            (tmr_registers(0)(429) and tmr_registers(2)(429));                                                         
                                                                                                                                     
        global_tmr_voter(0)(430)  <=    (tmr_registers(0)(430) and tmr_registers(1)(430)) or                                            
                            (tmr_registers(1)(430) and tmr_registers(2)(430)) or                                                       
                            (tmr_registers(0)(430) and tmr_registers(2)(430));                                                         
                                                                                                                                     
        global_tmr_voter(0)(431)  <=    (tmr_registers(0)(431) and tmr_registers(1)(431)) or                                            
                            (tmr_registers(1)(431) and tmr_registers(2)(431)) or                                                       
                            (tmr_registers(0)(431) and tmr_registers(2)(431));                                                         
                                                                                                                                     
        global_tmr_voter(0)(432)  <=    (tmr_registers(0)(432) and tmr_registers(1)(432)) or                                            
                            (tmr_registers(1)(432) and tmr_registers(2)(432)) or                                                       
                            (tmr_registers(0)(432) and tmr_registers(2)(432));                                                         
                                                                                                                                     
        global_tmr_voter(0)(433)  <=    (tmr_registers(0)(433) and tmr_registers(1)(433)) or                                            
                            (tmr_registers(1)(433) and tmr_registers(2)(433)) or                                                       
                            (tmr_registers(0)(433) and tmr_registers(2)(433));                                                         
                                                                                                                                     
        global_tmr_voter(0)(434)  <=    (tmr_registers(0)(434) and tmr_registers(1)(434)) or                                            
                            (tmr_registers(1)(434) and tmr_registers(2)(434)) or                                                       
                            (tmr_registers(0)(434) and tmr_registers(2)(434));                                                         
                                                                                                                                     
        global_tmr_voter(0)(435)  <=    (tmr_registers(0)(435) and tmr_registers(1)(435)) or                                            
                            (tmr_registers(1)(435) and tmr_registers(2)(435)) or                                                       
                            (tmr_registers(0)(435) and tmr_registers(2)(435));                                                         
                                                                                                                                     
        global_tmr_voter(0)(436)  <=    (tmr_registers(0)(436) and tmr_registers(1)(436)) or                                            
                            (tmr_registers(1)(436) and tmr_registers(2)(436)) or                                                       
                            (tmr_registers(0)(436) and tmr_registers(2)(436));                                                         
                                                                                                                                     
        global_tmr_voter(0)(437)  <=    (tmr_registers(0)(437) and tmr_registers(1)(437)) or                                            
                            (tmr_registers(1)(437) and tmr_registers(2)(437)) or                                                       
                            (tmr_registers(0)(437) and tmr_registers(2)(437));                                                         
                                                                                                                                     
        global_tmr_voter(0)(438)  <=    (tmr_registers(0)(438) and tmr_registers(1)(438)) or                                            
                            (tmr_registers(1)(438) and tmr_registers(2)(438)) or                                                       
                            (tmr_registers(0)(438) and tmr_registers(2)(438));                                                         
                                                                                                                                     
        global_tmr_voter(0)(439)  <=    (tmr_registers(0)(439) and tmr_registers(1)(439)) or                                            
                            (tmr_registers(1)(439) and tmr_registers(2)(439)) or                                                       
                            (tmr_registers(0)(439) and tmr_registers(2)(439));                                                         
                                                                                                                                     
        global_tmr_voter(0)(440)  <=    (tmr_registers(0)(440) and tmr_registers(1)(440)) or                                            
                            (tmr_registers(1)(440) and tmr_registers(2)(440)) or                                                       
                            (tmr_registers(0)(440) and tmr_registers(2)(440));                                                         
                                                                                                                                     
        global_tmr_voter(0)(441)  <=    (tmr_registers(0)(441) and tmr_registers(1)(441)) or                                            
                            (tmr_registers(1)(441) and tmr_registers(2)(441)) or                                                       
                            (tmr_registers(0)(441) and tmr_registers(2)(441));                                                         
                                                                                                                                     
        global_tmr_voter(0)(442)  <=    (tmr_registers(0)(442) and tmr_registers(1)(442)) or                                            
                            (tmr_registers(1)(442) and tmr_registers(2)(442)) or                                                       
                            (tmr_registers(0)(442) and tmr_registers(2)(442));                                                         
                                                                                                                                     
        global_tmr_voter(0)(443)  <=    (tmr_registers(0)(443) and tmr_registers(1)(443)) or                                            
                            (tmr_registers(1)(443) and tmr_registers(2)(443)) or                                                       
                            (tmr_registers(0)(443) and tmr_registers(2)(443));                                                         
                                                                                                                                     
        global_tmr_voter(0)(444)  <=    (tmr_registers(0)(444) and tmr_registers(1)(444)) or                                            
                            (tmr_registers(1)(444) and tmr_registers(2)(444)) or                                                       
                            (tmr_registers(0)(444) and tmr_registers(2)(444));                                                         
                                                                                                                                     
        global_tmr_voter(0)(445)  <=    (tmr_registers(0)(445) and tmr_registers(1)(445)) or                                            
                            (tmr_registers(1)(445) and tmr_registers(2)(445)) or                                                       
                            (tmr_registers(0)(445) and tmr_registers(2)(445));                                                         
                                                                                                                                     
        global_tmr_voter(0)(446)  <=    (tmr_registers(0)(446) and tmr_registers(1)(446)) or                                            
                            (tmr_registers(1)(446) and tmr_registers(2)(446)) or                                                       
                            (tmr_registers(0)(446) and tmr_registers(2)(446));                                                         
                                                                                                                                     
        global_tmr_voter(0)(447)  <=    (tmr_registers(0)(447) and tmr_registers(1)(447)) or                                            
                            (tmr_registers(1)(447) and tmr_registers(2)(447)) or                                                       
                            (tmr_registers(0)(447) and tmr_registers(2)(447));                                                         
                                                                                                                                     
        global_tmr_voter(0)(448)  <=    (tmr_registers(0)(448) and tmr_registers(1)(448)) or                                            
                            (tmr_registers(1)(448) and tmr_registers(2)(448)) or                                                       
                            (tmr_registers(0)(448) and tmr_registers(2)(448));                                                         
                                                                                                                                     
        global_tmr_voter(0)(449)  <=    (tmr_registers(0)(449) and tmr_registers(1)(449)) or                                            
                            (tmr_registers(1)(449) and tmr_registers(2)(449)) or                                                       
                            (tmr_registers(0)(449) and tmr_registers(2)(449));                                                         
                                                                                                                                     
        global_tmr_voter(0)(450)  <=    (tmr_registers(0)(450) and tmr_registers(1)(450)) or                                            
                            (tmr_registers(1)(450) and tmr_registers(2)(450)) or                                                       
                            (tmr_registers(0)(450) and tmr_registers(2)(450));                                                         
                                                                                                                                     
        global_tmr_voter(0)(451)  <=    (tmr_registers(0)(451) and tmr_registers(1)(451)) or                                            
                            (tmr_registers(1)(451) and tmr_registers(2)(451)) or                                                       
                            (tmr_registers(0)(451) and tmr_registers(2)(451));                                                         
                                                                                                                                     
        global_tmr_voter(0)(452)  <=    (tmr_registers(0)(452) and tmr_registers(1)(452)) or                                            
                            (tmr_registers(1)(452) and tmr_registers(2)(452)) or                                                       
                            (tmr_registers(0)(452) and tmr_registers(2)(452));                                                         
                                                                                                                                     
        global_tmr_voter(0)(453)  <=    (tmr_registers(0)(453) and tmr_registers(1)(453)) or                                            
                            (tmr_registers(1)(453) and tmr_registers(2)(453)) or                                                       
                            (tmr_registers(0)(453) and tmr_registers(2)(453));                                                         
                                                                                                                                     
        global_tmr_voter(0)(454)  <=    (tmr_registers(0)(454) and tmr_registers(1)(454)) or                                            
                            (tmr_registers(1)(454) and tmr_registers(2)(454)) or                                                       
                            (tmr_registers(0)(454) and tmr_registers(2)(454));                                                         
                                                                                                                                     
        global_tmr_voter(0)(455)  <=    (tmr_registers(0)(455) and tmr_registers(1)(455)) or                                            
                            (tmr_registers(1)(455) and tmr_registers(2)(455)) or                                                       
                            (tmr_registers(0)(455) and tmr_registers(2)(455));                                                         
                                                                                                                                     
        global_tmr_voter(0)(456)  <=    (tmr_registers(0)(456) and tmr_registers(1)(456)) or                                            
                            (tmr_registers(1)(456) and tmr_registers(2)(456)) or                                                       
                            (tmr_registers(0)(456) and tmr_registers(2)(456));                                                         
                                                                                                                                     
        global_tmr_voter(0)(457)  <=    (tmr_registers(0)(457) and tmr_registers(1)(457)) or                                            
                            (tmr_registers(1)(457) and tmr_registers(2)(457)) or                                                       
                            (tmr_registers(0)(457) and tmr_registers(2)(457));                                                         
                                                                                                                                     
        global_tmr_voter(0)(458)  <=    (tmr_registers(0)(458) and tmr_registers(1)(458)) or                                            
                            (tmr_registers(1)(458) and tmr_registers(2)(458)) or                                                       
                            (tmr_registers(0)(458) and tmr_registers(2)(458));                                                         
                                                                                                                                     
        global_tmr_voter(0)(459)  <=    (tmr_registers(0)(459) and tmr_registers(1)(459)) or                                            
                            (tmr_registers(1)(459) and tmr_registers(2)(459)) or                                                       
                            (tmr_registers(0)(459) and tmr_registers(2)(459));                                                         
                                                                                                                                     
        global_tmr_voter(0)(460)  <=    (tmr_registers(0)(460) and tmr_registers(1)(460)) or                                            
                            (tmr_registers(1)(460) and tmr_registers(2)(460)) or                                                       
                            (tmr_registers(0)(460) and tmr_registers(2)(460));                                                         
                                                                                                                                     
        global_tmr_voter(0)(461)  <=    (tmr_registers(0)(461) and tmr_registers(1)(461)) or                                            
                            (tmr_registers(1)(461) and tmr_registers(2)(461)) or                                                       
                            (tmr_registers(0)(461) and tmr_registers(2)(461));                                                         
                                                                                                                                     
        global_tmr_voter(0)(462)  <=    (tmr_registers(0)(462) and tmr_registers(1)(462)) or                                            
                            (tmr_registers(1)(462) and tmr_registers(2)(462)) or                                                       
                            (tmr_registers(0)(462) and tmr_registers(2)(462));                                                         
                                                                                                                                     
        global_tmr_voter(0)(463)  <=    (tmr_registers(0)(463) and tmr_registers(1)(463)) or                                            
                            (tmr_registers(1)(463) and tmr_registers(2)(463)) or                                                       
                            (tmr_registers(0)(463) and tmr_registers(2)(463));                                                         
                                                                                                                                     
        global_tmr_voter(0)(464)  <=    (tmr_registers(0)(464) and tmr_registers(1)(464)) or                                            
                            (tmr_registers(1)(464) and tmr_registers(2)(464)) or                                                       
                            (tmr_registers(0)(464) and tmr_registers(2)(464));                                                         
                                                                                                                                     
        global_tmr_voter(0)(465)  <=    (tmr_registers(0)(465) and tmr_registers(1)(465)) or                                            
                            (tmr_registers(1)(465) and tmr_registers(2)(465)) or                                                       
                            (tmr_registers(0)(465) and tmr_registers(2)(465));                                                         
                                                                                                                                     
        global_tmr_voter(0)(466)  <=    (tmr_registers(0)(466) and tmr_registers(1)(466)) or                                            
                            (tmr_registers(1)(466) and tmr_registers(2)(466)) or                                                       
                            (tmr_registers(0)(466) and tmr_registers(2)(466));                                                         
                                                                                                                                     
        global_tmr_voter(0)(467)  <=    (tmr_registers(0)(467) and tmr_registers(1)(467)) or                                            
                            (tmr_registers(1)(467) and tmr_registers(2)(467)) or                                                       
                            (tmr_registers(0)(467) and tmr_registers(2)(467));                                                         
                                                                                                                                     
        global_tmr_voter(0)(468)  <=    (tmr_registers(0)(468) and tmr_registers(1)(468)) or                                            
                            (tmr_registers(1)(468) and tmr_registers(2)(468)) or                                                       
                            (tmr_registers(0)(468) and tmr_registers(2)(468));                                                         
                                                                                                                                     
        global_tmr_voter(0)(469)  <=    (tmr_registers(0)(469) and tmr_registers(1)(469)) or                                            
                            (tmr_registers(1)(469) and tmr_registers(2)(469)) or                                                       
                            (tmr_registers(0)(469) and tmr_registers(2)(469));                                                         
                                                                                                                                     
        global_tmr_voter(0)(470)  <=    (tmr_registers(0)(470) and tmr_registers(1)(470)) or                                            
                            (tmr_registers(1)(470) and tmr_registers(2)(470)) or                                                       
                            (tmr_registers(0)(470) and tmr_registers(2)(470));                                                         
                                                                                                                                     
        global_tmr_voter(0)(471)  <=    (tmr_registers(0)(471) and tmr_registers(1)(471)) or                                            
                            (tmr_registers(1)(471) and tmr_registers(2)(471)) or                                                       
                            (tmr_registers(0)(471) and tmr_registers(2)(471));                                                         
                                                                                                                                     
        global_tmr_voter(0)(472)  <=    (tmr_registers(0)(472) and tmr_registers(1)(472)) or                                            
                            (tmr_registers(1)(472) and tmr_registers(2)(472)) or                                                       
                            (tmr_registers(0)(472) and tmr_registers(2)(472));                                                         
                                                                                                                                     
        global_tmr_voter(0)(473)  <=    (tmr_registers(0)(473) and tmr_registers(1)(473)) or                                            
                            (tmr_registers(1)(473) and tmr_registers(2)(473)) or                                                       
                            (tmr_registers(0)(473) and tmr_registers(2)(473));                                                         
                                                                                                                                     
        global_tmr_voter(0)(474)  <=    (tmr_registers(0)(474) and tmr_registers(1)(474)) or                                            
                            (tmr_registers(1)(474) and tmr_registers(2)(474)) or                                                       
                            (tmr_registers(0)(474) and tmr_registers(2)(474));                                                         
                                                                                                                                     
        global_tmr_voter(0)(475)  <=    (tmr_registers(0)(475) and tmr_registers(1)(475)) or                                            
                            (tmr_registers(1)(475) and tmr_registers(2)(475)) or                                                       
                            (tmr_registers(0)(475) and tmr_registers(2)(475));                                                         
                                                                                                                                     
        global_tmr_voter(0)(476)  <=    (tmr_registers(0)(476) and tmr_registers(1)(476)) or                                            
                            (tmr_registers(1)(476) and tmr_registers(2)(476)) or                                                       
                            (tmr_registers(0)(476) and tmr_registers(2)(476));                                                         
                                                                                                                                     
        global_tmr_voter(0)(477)  <=    (tmr_registers(0)(477) and tmr_registers(1)(477)) or                                            
                            (tmr_registers(1)(477) and tmr_registers(2)(477)) or                                                       
                            (tmr_registers(0)(477) and tmr_registers(2)(477));                                                         
                                                                                                                                     
        global_tmr_voter(0)(478)  <=    (tmr_registers(0)(478) and tmr_registers(1)(478)) or                                            
                            (tmr_registers(1)(478) and tmr_registers(2)(478)) or                                                       
                            (tmr_registers(0)(478) and tmr_registers(2)(478));                                                         
                                                                                                                                     
        global_tmr_voter(0)(479)  <=    (tmr_registers(0)(479) and tmr_registers(1)(479)) or                                            
                            (tmr_registers(1)(479) and tmr_registers(2)(479)) or                                                       
                            (tmr_registers(0)(479) and tmr_registers(2)(479));                                                         
                                                                                                                                     
        global_tmr_voter(0)(480)  <=    (tmr_registers(0)(480) and tmr_registers(1)(480)) or                                            
                            (tmr_registers(1)(480) and tmr_registers(2)(480)) or                                                       
                            (tmr_registers(0)(480) and tmr_registers(2)(480));                                                         
                                                                                                                                     
        global_tmr_voter(0)(481)  <=    (tmr_registers(0)(481) and tmr_registers(1)(481)) or                                            
                            (tmr_registers(1)(481) and tmr_registers(2)(481)) or                                                       
                            (tmr_registers(0)(481) and tmr_registers(2)(481));                                                         
                                                                                                                                     
        global_tmr_voter(0)(482)  <=    (tmr_registers(0)(482) and tmr_registers(1)(482)) or                                            
                            (tmr_registers(1)(482) and tmr_registers(2)(482)) or                                                       
                            (tmr_registers(0)(482) and tmr_registers(2)(482));                                                         
                                                                                                                                     
        global_tmr_voter(0)(483)  <=    (tmr_registers(0)(483) and tmr_registers(1)(483)) or                                            
                            (tmr_registers(1)(483) and tmr_registers(2)(483)) or                                                       
                            (tmr_registers(0)(483) and tmr_registers(2)(483));                                                         
                                                                                                                                     
        global_tmr_voter(0)(484)  <=    (tmr_registers(0)(484) and tmr_registers(1)(484)) or                                            
                            (tmr_registers(1)(484) and tmr_registers(2)(484)) or                                                       
                            (tmr_registers(0)(484) and tmr_registers(2)(484));                                                         
                                                                                                                                     
        global_tmr_voter(0)(485)  <=    (tmr_registers(0)(485) and tmr_registers(1)(485)) or                                            
                            (tmr_registers(1)(485) and tmr_registers(2)(485)) or                                                       
                            (tmr_registers(0)(485) and tmr_registers(2)(485));                                                         
                                                                                                                                     
        global_tmr_voter(0)(486)  <=    (tmr_registers(0)(486) and tmr_registers(1)(486)) or                                            
                            (tmr_registers(1)(486) and tmr_registers(2)(486)) or                                                       
                            (tmr_registers(0)(486) and tmr_registers(2)(486));                                                         
                                                                                                                                     
        global_tmr_voter(0)(487)  <=    (tmr_registers(0)(487) and tmr_registers(1)(487)) or                                            
                            (tmr_registers(1)(487) and tmr_registers(2)(487)) or                                                       
                            (tmr_registers(0)(487) and tmr_registers(2)(487));                                                         
                                                                                                                                     
        global_tmr_voter(0)(488)  <=    (tmr_registers(0)(488) and tmr_registers(1)(488)) or                                            
                            (tmr_registers(1)(488) and tmr_registers(2)(488)) or                                                       
                            (tmr_registers(0)(488) and tmr_registers(2)(488));                                                         
                                                                                                                                     
        global_tmr_voter(0)(489)  <=    (tmr_registers(0)(489) and tmr_registers(1)(489)) or                                            
                            (tmr_registers(1)(489) and tmr_registers(2)(489)) or                                                       
                            (tmr_registers(0)(489) and tmr_registers(2)(489));                                                         
                                                                                                                                     
        global_tmr_voter(0)(490)  <=    (tmr_registers(0)(490) and tmr_registers(1)(490)) or                                            
                            (tmr_registers(1)(490) and tmr_registers(2)(490)) or                                                       
                            (tmr_registers(0)(490) and tmr_registers(2)(490));                                                         
                                                                                                                                     
        global_tmr_voter(0)(491)  <=    (tmr_registers(0)(491) and tmr_registers(1)(491)) or                                            
                            (tmr_registers(1)(491) and tmr_registers(2)(491)) or                                                       
                            (tmr_registers(0)(491) and tmr_registers(2)(491));                                                         
                                                                                                                                     
        global_tmr_voter(0)(492)  <=    (tmr_registers(0)(492) and tmr_registers(1)(492)) or                                            
                            (tmr_registers(1)(492) and tmr_registers(2)(492)) or                                                       
                            (tmr_registers(0)(492) and tmr_registers(2)(492));                                                         
                                                                                                                                     
        global_tmr_voter(0)(493)  <=    (tmr_registers(0)(493) and tmr_registers(1)(493)) or                                            
                            (tmr_registers(1)(493) and tmr_registers(2)(493)) or                                                       
                            (tmr_registers(0)(493) and tmr_registers(2)(493));                                                         
                                                                                                                                     
        global_tmr_voter(0)(494)  <=    (tmr_registers(0)(494) and tmr_registers(1)(494)) or                                            
                            (tmr_registers(1)(494) and tmr_registers(2)(494)) or                                                       
                            (tmr_registers(0)(494) and tmr_registers(2)(494));                                                         
                                                                                                                                     
        global_tmr_voter(0)(495)  <=    (tmr_registers(0)(495) and tmr_registers(1)(495)) or                                            
                            (tmr_registers(1)(495) and tmr_registers(2)(495)) or                                                       
                            (tmr_registers(0)(495) and tmr_registers(2)(495));                                                         
                                                                                                                                     
        global_tmr_voter(0)(496)  <=    (tmr_registers(0)(496) and tmr_registers(1)(496)) or                                            
                            (tmr_registers(1)(496) and tmr_registers(2)(496)) or                                                       
                            (tmr_registers(0)(496) and tmr_registers(2)(496));                                                         
                                                                                                                                     
        global_tmr_voter(0)(497)  <=    (tmr_registers(0)(497) and tmr_registers(1)(497)) or                                            
                            (tmr_registers(1)(497) and tmr_registers(2)(497)) or                                                       
                            (tmr_registers(0)(497) and tmr_registers(2)(497));                                                         
                                                                                                                                     
        global_tmr_voter(0)(498)  <=    (tmr_registers(0)(498) and tmr_registers(1)(498)) or                                            
                            (tmr_registers(1)(498) and tmr_registers(2)(498)) or                                                       
                            (tmr_registers(0)(498) and tmr_registers(2)(498));                                                         
                                                                                                                                     
        global_tmr_voter(0)(499)  <=    (tmr_registers(0)(499) and tmr_registers(1)(499)) or                                            
                            (tmr_registers(1)(499) and tmr_registers(2)(499)) or                                                       
                            (tmr_registers(0)(499) and tmr_registers(2)(499));                                                         
                                                                                                                                     
        global_tmr_voter(0)(500)  <=    (tmr_registers(0)(500) and tmr_registers(1)(500)) or                                            
                            (tmr_registers(1)(500) and tmr_registers(2)(500)) or                                                       
                            (tmr_registers(0)(500) and tmr_registers(2)(500));                                                         
                                                                                                                                     
        global_tmr_voter(0)(501)  <=    (tmr_registers(0)(501) and tmr_registers(1)(501)) or                                            
                            (tmr_registers(1)(501) and tmr_registers(2)(501)) or                                                       
                            (tmr_registers(0)(501) and tmr_registers(2)(501));                                                         
                                                                                                                                     
        global_tmr_voter(0)(502)  <=    (tmr_registers(0)(502) and tmr_registers(1)(502)) or                                            
                            (tmr_registers(1)(502) and tmr_registers(2)(502)) or                                                       
                            (tmr_registers(0)(502) and tmr_registers(2)(502));                                                         
                                                                                                                                     
        global_tmr_voter(0)(503)  <=    (tmr_registers(0)(503) and tmr_registers(1)(503)) or                                            
                            (tmr_registers(1)(503) and tmr_registers(2)(503)) or                                                       
                            (tmr_registers(0)(503) and tmr_registers(2)(503));                                                         
                                                                                                                                     
        global_tmr_voter(0)(504)  <=    (tmr_registers(0)(504) and tmr_registers(1)(504)) or                                            
                            (tmr_registers(1)(504) and tmr_registers(2)(504)) or                                                       
                            (tmr_registers(0)(504) and tmr_registers(2)(504));                                                         
                                                                                                                                     
        global_tmr_voter(0)(505)  <=    (tmr_registers(0)(505) and tmr_registers(1)(505)) or                                            
                            (tmr_registers(1)(505) and tmr_registers(2)(505)) or                                                       
                            (tmr_registers(0)(505) and tmr_registers(2)(505));                                                         
                                                                                                                                     
        global_tmr_voter(0)(506)  <=    (tmr_registers(0)(506) and tmr_registers(1)(506)) or                                            
                            (tmr_registers(1)(506) and tmr_registers(2)(506)) or                                                       
                            (tmr_registers(0)(506) and tmr_registers(2)(506));                                                         
                                                                                                                                     
        global_tmr_voter(0)(507)  <=    (tmr_registers(0)(507) and tmr_registers(1)(507)) or                                            
                            (tmr_registers(1)(507) and tmr_registers(2)(507)) or                                                       
                            (tmr_registers(0)(507) and tmr_registers(2)(507));                                                         
                                                                                                                                     
        global_tmr_voter(0)(508)  <=    (tmr_registers(0)(508) and tmr_registers(1)(508)) or                                            
                            (tmr_registers(1)(508) and tmr_registers(2)(508)) or                                                       
                            (tmr_registers(0)(508) and tmr_registers(2)(508));                                                         
                                                                                                                                     
        global_tmr_voter(0)(509)  <=    (tmr_registers(0)(509) and tmr_registers(1)(509)) or                                            
                            (tmr_registers(1)(509) and tmr_registers(2)(509)) or                                                       
                            (tmr_registers(0)(509) and tmr_registers(2)(509));                                                         
                                                                                                                                     
        global_tmr_voter(0)(510)  <=    (tmr_registers(0)(510) and tmr_registers(1)(510)) or                                            
                            (tmr_registers(1)(510) and tmr_registers(2)(510)) or                                                       
                            (tmr_registers(0)(510) and tmr_registers(2)(510));                                                         
                                                                                                                                     
        global_tmr_voter(0)(511)  <=    (tmr_registers(0)(511) and tmr_registers(1)(511)) or                                            
                            (tmr_registers(1)(511) and tmr_registers(2)(511)) or                                                       
                            (tmr_registers(0)(511) and tmr_registers(2)(511));                                                         
                                                                                                                                     
        global_tmr_voter(0)(512)  <=    (tmr_registers(0)(512) and tmr_registers(1)(512)) or                                            
                            (tmr_registers(1)(512) and tmr_registers(2)(512)) or                                                       
                            (tmr_registers(0)(512) and tmr_registers(2)(512));                                                         
                                                                                                                                     
        global_tmr_voter(0)(513)  <=    (tmr_registers(0)(513) and tmr_registers(1)(513)) or                                            
                            (tmr_registers(1)(513) and tmr_registers(2)(513)) or                                                       
                            (tmr_registers(0)(513) and tmr_registers(2)(513));                                                         
                                                                                                                                     
        global_tmr_voter(0)(514)  <=    (tmr_registers(0)(514) and tmr_registers(1)(514)) or                                            
                            (tmr_registers(1)(514) and tmr_registers(2)(514)) or                                                       
                            (tmr_registers(0)(514) and tmr_registers(2)(514));                                                         
                                                                                                                                     
        global_tmr_voter(0)(515)  <=    (tmr_registers(0)(515) and tmr_registers(1)(515)) or                                            
                            (tmr_registers(1)(515) and tmr_registers(2)(515)) or                                                       
                            (tmr_registers(0)(515) and tmr_registers(2)(515));                                                         
                                                                                                                                     
        global_tmr_voter(0)(516)  <=    (tmr_registers(0)(516) and tmr_registers(1)(516)) or                                            
                            (tmr_registers(1)(516) and tmr_registers(2)(516)) or                                                       
                            (tmr_registers(0)(516) and tmr_registers(2)(516));                                                         
                                                                                                                                     
        global_tmr_voter(0)(517)  <=    (tmr_registers(0)(517) and tmr_registers(1)(517)) or                                            
                            (tmr_registers(1)(517) and tmr_registers(2)(517)) or                                                       
                            (tmr_registers(0)(517) and tmr_registers(2)(517));                                                         
                                                                                                                                     
        global_tmr_voter(0)(518)  <=    (tmr_registers(0)(518) and tmr_registers(1)(518)) or                                            
                            (tmr_registers(1)(518) and tmr_registers(2)(518)) or                                                       
                            (tmr_registers(0)(518) and tmr_registers(2)(518));                                                         
                                                                                                                                     
        global_tmr_voter(0)(519)  <=    (tmr_registers(0)(519) and tmr_registers(1)(519)) or                                            
                            (tmr_registers(1)(519) and tmr_registers(2)(519)) or                                                       
                            (tmr_registers(0)(519) and tmr_registers(2)(519));                                                         
                                                                                                                                     
        global_tmr_voter(0)(520)  <=    (tmr_registers(0)(520) and tmr_registers(1)(520)) or                                            
                            (tmr_registers(1)(520) and tmr_registers(2)(520)) or                                                       
                            (tmr_registers(0)(520) and tmr_registers(2)(520));                                                         
                                                                                                                                     
        global_tmr_voter(0)(521)  <=    (tmr_registers(0)(521) and tmr_registers(1)(521)) or                                            
                            (tmr_registers(1)(521) and tmr_registers(2)(521)) or                                                       
                            (tmr_registers(0)(521) and tmr_registers(2)(521));                                                         
                                                                                                                                     
        global_tmr_voter(0)(522)  <=    (tmr_registers(0)(522) and tmr_registers(1)(522)) or                                            
                            (tmr_registers(1)(522) and tmr_registers(2)(522)) or                                                       
                            (tmr_registers(0)(522) and tmr_registers(2)(522));                                                         
                                                                                                                                     
        global_tmr_voter(0)(523)  <=    (tmr_registers(0)(523) and tmr_registers(1)(523)) or                                            
                            (tmr_registers(1)(523) and tmr_registers(2)(523)) or                                                       
                            (tmr_registers(0)(523) and tmr_registers(2)(523));                                                         
                                                                                                                                     
        global_tmr_voter(0)(524)  <=    (tmr_registers(0)(524) and tmr_registers(1)(524)) or                                            
                            (tmr_registers(1)(524) and tmr_registers(2)(524)) or                                                       
                            (tmr_registers(0)(524) and tmr_registers(2)(524));                                                         
                                                                                                                                     
        global_tmr_voter(0)(525)  <=    (tmr_registers(0)(525) and tmr_registers(1)(525)) or                                            
                            (tmr_registers(1)(525) and tmr_registers(2)(525)) or                                                       
                            (tmr_registers(0)(525) and tmr_registers(2)(525));                                                         
                                                                                                                                     
        global_tmr_voter(0)(526)  <=    (tmr_registers(0)(526) and tmr_registers(1)(526)) or                                            
                            (tmr_registers(1)(526) and tmr_registers(2)(526)) or                                                       
                            (tmr_registers(0)(526) and tmr_registers(2)(526));                                                         
                                                                                                                                     
        global_tmr_voter(0)(527)  <=    (tmr_registers(0)(527) and tmr_registers(1)(527)) or                                            
                            (tmr_registers(1)(527) and tmr_registers(2)(527)) or                                                       
                            (tmr_registers(0)(527) and tmr_registers(2)(527));                                                         
                                                                                                                                     
        global_tmr_voter(0)(528)  <=    (tmr_registers(0)(528) and tmr_registers(1)(528)) or                                            
                            (tmr_registers(1)(528) and tmr_registers(2)(528)) or                                                       
                            (tmr_registers(0)(528) and tmr_registers(2)(528));                                                         
                                                                                                                                     
        global_tmr_voter(0)(529)  <=    (tmr_registers(0)(529) and tmr_registers(1)(529)) or                                            
                            (tmr_registers(1)(529) and tmr_registers(2)(529)) or                                                       
                            (tmr_registers(0)(529) and tmr_registers(2)(529));                                                         
                                                                                                                                     
        global_tmr_voter(0)(530)  <=    (tmr_registers(0)(530) and tmr_registers(1)(530)) or                                            
                            (tmr_registers(1)(530) and tmr_registers(2)(530)) or                                                       
                            (tmr_registers(0)(530) and tmr_registers(2)(530));                                                         
                                                                                                                                     
        global_tmr_voter(0)(531)  <=    (tmr_registers(0)(531) and tmr_registers(1)(531)) or                                            
                            (tmr_registers(1)(531) and tmr_registers(2)(531)) or                                                       
                            (tmr_registers(0)(531) and tmr_registers(2)(531));                                                         
                                                                                                                                     
        global_tmr_voter(0)(532)  <=    (tmr_registers(0)(532) and tmr_registers(1)(532)) or                                            
                            (tmr_registers(1)(532) and tmr_registers(2)(532)) or                                                       
                            (tmr_registers(0)(532) and tmr_registers(2)(532));                                                         
                                                                                                                                     
        global_tmr_voter(0)(533)  <=    (tmr_registers(0)(533) and tmr_registers(1)(533)) or                                            
                            (tmr_registers(1)(533) and tmr_registers(2)(533)) or                                                       
                            (tmr_registers(0)(533) and tmr_registers(2)(533));                                                         
                                                                                                                                     
        global_tmr_voter(0)(534)  <=    (tmr_registers(0)(534) and tmr_registers(1)(534)) or                                            
                            (tmr_registers(1)(534) and tmr_registers(2)(534)) or                                                       
                            (tmr_registers(0)(534) and tmr_registers(2)(534));                                                         
                                                                                                                                     
        global_tmr_voter(0)(535)  <=    (tmr_registers(0)(535) and tmr_registers(1)(535)) or                                            
                            (tmr_registers(1)(535) and tmr_registers(2)(535)) or                                                       
                            (tmr_registers(0)(535) and tmr_registers(2)(535));                                                         
                                                                                                                                     
        global_tmr_voter(0)(536)  <=    (tmr_registers(0)(536) and tmr_registers(1)(536)) or                                            
                            (tmr_registers(1)(536) and tmr_registers(2)(536)) or                                                       
                            (tmr_registers(0)(536) and tmr_registers(2)(536));                                                         
                                                                                                                                     
        global_tmr_voter(0)(537)  <=    (tmr_registers(0)(537) and tmr_registers(1)(537)) or                                            
                            (tmr_registers(1)(537) and tmr_registers(2)(537)) or                                                       
                            (tmr_registers(0)(537) and tmr_registers(2)(537));                                                         
                                                                                                                                     
        global_tmr_voter(0)(538)  <=    (tmr_registers(0)(538) and tmr_registers(1)(538)) or                                            
                            (tmr_registers(1)(538) and tmr_registers(2)(538)) or                                                       
                            (tmr_registers(0)(538) and tmr_registers(2)(538));                                                         
                                                                                                                                     
        global_tmr_voter(0)(539)  <=    (tmr_registers(0)(539) and tmr_registers(1)(539)) or                                            
                            (tmr_registers(1)(539) and tmr_registers(2)(539)) or                                                       
                            (tmr_registers(0)(539) and tmr_registers(2)(539));                                                         
                                                                                                                                     
        global_tmr_voter(0)(540)  <=    (tmr_registers(0)(540) and tmr_registers(1)(540)) or                                            
                            (tmr_registers(1)(540) and tmr_registers(2)(540)) or                                                       
                            (tmr_registers(0)(540) and tmr_registers(2)(540));                                                         
                                                                                                                                     
        global_tmr_voter(0)(541)  <=    (tmr_registers(0)(541) and tmr_registers(1)(541)) or                                            
                            (tmr_registers(1)(541) and tmr_registers(2)(541)) or                                                       
                            (tmr_registers(0)(541) and tmr_registers(2)(541));                                                         
                                                                                                                                     
        global_tmr_voter(0)(542)  <=    (tmr_registers(0)(542) and tmr_registers(1)(542)) or                                            
                            (tmr_registers(1)(542) and tmr_registers(2)(542)) or                                                       
                            (tmr_registers(0)(542) and tmr_registers(2)(542));                                                         
                                                                                                                                     
        global_tmr_voter(0)(543)  <=    (tmr_registers(0)(543) and tmr_registers(1)(543)) or                                            
                            (tmr_registers(1)(543) and tmr_registers(2)(543)) or                                                       
                            (tmr_registers(0)(543) and tmr_registers(2)(543));                                                         
                                                                                                                                     
        global_tmr_voter(0)(544)  <=    (tmr_registers(0)(544) and tmr_registers(1)(544)) or                                            
                            (tmr_registers(1)(544) and tmr_registers(2)(544)) or                                                       
                            (tmr_registers(0)(544) and tmr_registers(2)(544));                                                         
                                                                                                                                     
        global_tmr_voter(0)(545)  <=    (tmr_registers(0)(545) and tmr_registers(1)(545)) or                                            
                            (tmr_registers(1)(545) and tmr_registers(2)(545)) or                                                       
                            (tmr_registers(0)(545) and tmr_registers(2)(545));                                                         
                                                                                                                                     
        global_tmr_voter(0)(546)  <=    (tmr_registers(0)(546) and tmr_registers(1)(546)) or                                            
                            (tmr_registers(1)(546) and tmr_registers(2)(546)) or                                                       
                            (tmr_registers(0)(546) and tmr_registers(2)(546));                                                         
                                                                                                                                     
        global_tmr_voter(0)(547)  <=    (tmr_registers(0)(547) and tmr_registers(1)(547)) or                                            
                            (tmr_registers(1)(547) and tmr_registers(2)(547)) or                                                       
                            (tmr_registers(0)(547) and tmr_registers(2)(547));                                                         
                                                                                                                                     
        global_tmr_voter(0)(548)  <=    (tmr_registers(0)(548) and tmr_registers(1)(548)) or                                            
                            (tmr_registers(1)(548) and tmr_registers(2)(548)) or                                                       
                            (tmr_registers(0)(548) and tmr_registers(2)(548));                                                         
                                                                                                                                     
        global_tmr_voter(0)(549)  <=    (tmr_registers(0)(549) and tmr_registers(1)(549)) or                                            
                            (tmr_registers(1)(549) and tmr_registers(2)(549)) or                                                       
                            (tmr_registers(0)(549) and tmr_registers(2)(549));                                                         
                                                                                                                                     
        global_tmr_voter(0)(550)  <=    (tmr_registers(0)(550) and tmr_registers(1)(550)) or                                            
                            (tmr_registers(1)(550) and tmr_registers(2)(550)) or                                                       
                            (tmr_registers(0)(550) and tmr_registers(2)(550));                                                         
                                                                                                                                     
        global_tmr_voter(0)(551)  <=    (tmr_registers(0)(551) and tmr_registers(1)(551)) or                                            
                            (tmr_registers(1)(551) and tmr_registers(2)(551)) or                                                       
                            (tmr_registers(0)(551) and tmr_registers(2)(551));                                                         
                                                                                                                                     
        global_tmr_voter(0)(552)  <=    (tmr_registers(0)(552) and tmr_registers(1)(552)) or                                            
                            (tmr_registers(1)(552) and tmr_registers(2)(552)) or                                                       
                            (tmr_registers(0)(552) and tmr_registers(2)(552));                                                         
                                                                                                                                     
        global_tmr_voter(0)(553)  <=    (tmr_registers(0)(553) and tmr_registers(1)(553)) or                                            
                            (tmr_registers(1)(553) and tmr_registers(2)(553)) or                                                       
                            (tmr_registers(0)(553) and tmr_registers(2)(553));                                                         
                                                                                                                                     
        global_tmr_voter(0)(554)  <=    (tmr_registers(0)(554) and tmr_registers(1)(554)) or                                            
                            (tmr_registers(1)(554) and tmr_registers(2)(554)) or                                                       
                            (tmr_registers(0)(554) and tmr_registers(2)(554));                                                         
                                                                                                                                     
        global_tmr_voter(0)(555)  <=    (tmr_registers(0)(555) and tmr_registers(1)(555)) or                                            
                            (tmr_registers(1)(555) and tmr_registers(2)(555)) or                                                       
                            (tmr_registers(0)(555) and tmr_registers(2)(555));                                                         
                                                                                                                                     
        global_tmr_voter(0)(556)  <=    (tmr_registers(0)(556) and tmr_registers(1)(556)) or                                            
                            (tmr_registers(1)(556) and tmr_registers(2)(556)) or                                                       
                            (tmr_registers(0)(556) and tmr_registers(2)(556));                                                         
                                                                                                                                     
        global_tmr_voter(0)(557)  <=    (tmr_registers(0)(557) and tmr_registers(1)(557)) or                                            
                            (tmr_registers(1)(557) and tmr_registers(2)(557)) or                                                       
                            (tmr_registers(0)(557) and tmr_registers(2)(557));                                                         
                                                                                                                                     
        global_tmr_voter(0)(558)  <=    (tmr_registers(0)(558) and tmr_registers(1)(558)) or                                            
                            (tmr_registers(1)(558) and tmr_registers(2)(558)) or                                                       
                            (tmr_registers(0)(558) and tmr_registers(2)(558));                                                         
                                                                                                                                     
        global_tmr_voter(0)(559)  <=    (tmr_registers(0)(559) and tmr_registers(1)(559)) or                                            
                            (tmr_registers(1)(559) and tmr_registers(2)(559)) or                                                       
                            (tmr_registers(0)(559) and tmr_registers(2)(559));                                                         
                                                                                                                                     
        global_tmr_voter(0)(560)  <=    (tmr_registers(0)(560) and tmr_registers(1)(560)) or                                            
                            (tmr_registers(1)(560) and tmr_registers(2)(560)) or                                                       
                            (tmr_registers(0)(560) and tmr_registers(2)(560));                                                         
                                                                                                                                     
        global_tmr_voter(0)(561)  <=    (tmr_registers(0)(561) and tmr_registers(1)(561)) or                                            
                            (tmr_registers(1)(561) and tmr_registers(2)(561)) or                                                       
                            (tmr_registers(0)(561) and tmr_registers(2)(561));                                                         
                                                                                                                                     
        global_tmr_voter(0)(562)  <=    (tmr_registers(0)(562) and tmr_registers(1)(562)) or                                            
                            (tmr_registers(1)(562) and tmr_registers(2)(562)) or                                                       
                            (tmr_registers(0)(562) and tmr_registers(2)(562));                                                         
                                                                                                                                     
        global_tmr_voter(0)(563)  <=    (tmr_registers(0)(563) and tmr_registers(1)(563)) or                                            
                            (tmr_registers(1)(563) and tmr_registers(2)(563)) or                                                       
                            (tmr_registers(0)(563) and tmr_registers(2)(563));                                                         
                                                                                                                                     
        global_tmr_voter(0)(564)  <=    (tmr_registers(0)(564) and tmr_registers(1)(564)) or                                            
                            (tmr_registers(1)(564) and tmr_registers(2)(564)) or                                                       
                            (tmr_registers(0)(564) and tmr_registers(2)(564));                                                         
                                                                                                                                     
        global_tmr_voter(0)(565)  <=    (tmr_registers(0)(565) and tmr_registers(1)(565)) or                                            
                            (tmr_registers(1)(565) and tmr_registers(2)(565)) or                                                       
                            (tmr_registers(0)(565) and tmr_registers(2)(565));                                                         
                                                                                                                                     
        global_tmr_voter(0)(566)  <=    (tmr_registers(0)(566) and tmr_registers(1)(566)) or                                            
                            (tmr_registers(1)(566) and tmr_registers(2)(566)) or                                                       
                            (tmr_registers(0)(566) and tmr_registers(2)(566));                                                         
                                                                                                                                     
        global_tmr_voter(0)(567)  <=    (tmr_registers(0)(567) and tmr_registers(1)(567)) or                                            
                            (tmr_registers(1)(567) and tmr_registers(2)(567)) or                                                       
                            (tmr_registers(0)(567) and tmr_registers(2)(567));                                                         
                                                                                                                                     
        global_tmr_voter(0)(568)  <=    (tmr_registers(0)(568) and tmr_registers(1)(568)) or                                            
                            (tmr_registers(1)(568) and tmr_registers(2)(568)) or                                                       
                            (tmr_registers(0)(568) and tmr_registers(2)(568));                                                         
                                                                                                                                     
        global_tmr_voter(0)(569)  <=    (tmr_registers(0)(569) and tmr_registers(1)(569)) or                                            
                            (tmr_registers(1)(569) and tmr_registers(2)(569)) or                                                       
                            (tmr_registers(0)(569) and tmr_registers(2)(569));                                                         
                                                                                                                                     
        global_tmr_voter(0)(570)  <=    (tmr_registers(0)(570) and tmr_registers(1)(570)) or                                            
                            (tmr_registers(1)(570) and tmr_registers(2)(570)) or                                                       
                            (tmr_registers(0)(570) and tmr_registers(2)(570));                                                         
                                                                                                                                     
        global_tmr_voter(0)(571)  <=    (tmr_registers(0)(571) and tmr_registers(1)(571)) or                                            
                            (tmr_registers(1)(571) and tmr_registers(2)(571)) or                                                       
                            (tmr_registers(0)(571) and tmr_registers(2)(571));                                                         
                                                                                                                                     
        global_tmr_voter(0)(572)  <=    (tmr_registers(0)(572) and tmr_registers(1)(572)) or                                            
                            (tmr_registers(1)(572) and tmr_registers(2)(572)) or                                                       
                            (tmr_registers(0)(572) and tmr_registers(2)(572));                                                         
                                                                                                                                     
        global_tmr_voter(0)(573)  <=    (tmr_registers(0)(573) and tmr_registers(1)(573)) or                                            
                            (tmr_registers(1)(573) and tmr_registers(2)(573)) or                                                       
                            (tmr_registers(0)(573) and tmr_registers(2)(573));                                                         
                                                                                                                                     
        global_tmr_voter(0)(574)  <=    (tmr_registers(0)(574) and tmr_registers(1)(574)) or                                            
                            (tmr_registers(1)(574) and tmr_registers(2)(574)) or                                                       
                            (tmr_registers(0)(574) and tmr_registers(2)(574));                                                         
                                                                                                                                     
        global_tmr_voter(0)(575)  <=    (tmr_registers(0)(575) and tmr_registers(1)(575)) or                                            
                            (tmr_registers(1)(575) and tmr_registers(2)(575)) or                                                       
                            (tmr_registers(0)(575) and tmr_registers(2)(575));                                                         
                                                                                                                                     
        global_tmr_voter(0)(576)  <=    (tmr_registers(0)(576) and tmr_registers(1)(576)) or                                            
                            (tmr_registers(1)(576) and tmr_registers(2)(576)) or                                                       
                            (tmr_registers(0)(576) and tmr_registers(2)(576));                                                         
                                                                                                                                     
        global_tmr_voter(0)(577)  <=    (tmr_registers(0)(577) and tmr_registers(1)(577)) or                                            
                            (tmr_registers(1)(577) and tmr_registers(2)(577)) or                                                       
                            (tmr_registers(0)(577) and tmr_registers(2)(577));                                                         
                                                                                                                                     
        global_tmr_voter(0)(578)  <=    (tmr_registers(0)(578) and tmr_registers(1)(578)) or                                            
                            (tmr_registers(1)(578) and tmr_registers(2)(578)) or                                                       
                            (tmr_registers(0)(578) and tmr_registers(2)(578));                                                         
                                                                                                                                     
        global_tmr_voter(0)(579)  <=    (tmr_registers(0)(579) and tmr_registers(1)(579)) or                                            
                            (tmr_registers(1)(579) and tmr_registers(2)(579)) or                                                       
                            (tmr_registers(0)(579) and tmr_registers(2)(579));                                                         
                                                                                                                                     
        global_tmr_voter(0)(580)  <=    (tmr_registers(0)(580) and tmr_registers(1)(580)) or                                            
                            (tmr_registers(1)(580) and tmr_registers(2)(580)) or                                                       
                            (tmr_registers(0)(580) and tmr_registers(2)(580));                                                         
                                                                                                                                     
        global_tmr_voter(0)(581)  <=    (tmr_registers(0)(581) and tmr_registers(1)(581)) or                                            
                            (tmr_registers(1)(581) and tmr_registers(2)(581)) or                                                       
                            (tmr_registers(0)(581) and tmr_registers(2)(581));                                                         
                                                                                                                                     
        global_tmr_voter(0)(582)  <=    (tmr_registers(0)(582) and tmr_registers(1)(582)) or                                            
                            (tmr_registers(1)(582) and tmr_registers(2)(582)) or                                                       
                            (tmr_registers(0)(582) and tmr_registers(2)(582));                                                         
                                                                                                                                     
        global_tmr_voter(0)(583)  <=    (tmr_registers(0)(583) and tmr_registers(1)(583)) or                                            
                            (tmr_registers(1)(583) and tmr_registers(2)(583)) or                                                       
                            (tmr_registers(0)(583) and tmr_registers(2)(583));                                                         
                                                                                                                                     
        global_tmr_voter(0)(584)  <=    (tmr_registers(0)(584) and tmr_registers(1)(584)) or                                            
                            (tmr_registers(1)(584) and tmr_registers(2)(584)) or                                                       
                            (tmr_registers(0)(584) and tmr_registers(2)(584));                                                         
                                                                                                                                     
        global_tmr_voter(0)(585)  <=    (tmr_registers(0)(585) and tmr_registers(1)(585)) or                                            
                            (tmr_registers(1)(585) and tmr_registers(2)(585)) or                                                       
                            (tmr_registers(0)(585) and tmr_registers(2)(585));                                                         
                                                                                                                                     
        global_tmr_voter(0)(586)  <=    (tmr_registers(0)(586) and tmr_registers(1)(586)) or                                            
                            (tmr_registers(1)(586) and tmr_registers(2)(586)) or                                                       
                            (tmr_registers(0)(586) and tmr_registers(2)(586));                                                         
                                                                                                                                     
        global_tmr_voter(0)(587)  <=    (tmr_registers(0)(587) and tmr_registers(1)(587)) or                                            
                            (tmr_registers(1)(587) and tmr_registers(2)(587)) or                                                       
                            (tmr_registers(0)(587) and tmr_registers(2)(587));                                                         
                                                                                                                                     
        global_tmr_voter(0)(588)  <=    (tmr_registers(0)(588) and tmr_registers(1)(588)) or                                            
                            (tmr_registers(1)(588) and tmr_registers(2)(588)) or                                                       
                            (tmr_registers(0)(588) and tmr_registers(2)(588));                                                         
                                                                                                                                     
        global_tmr_voter(0)(589)  <=    (tmr_registers(0)(589) and tmr_registers(1)(589)) or                                            
                            (tmr_registers(1)(589) and tmr_registers(2)(589)) or                                                       
                            (tmr_registers(0)(589) and tmr_registers(2)(589));                                                         
                                                                                                                                     
        global_tmr_voter(0)(590)  <=    (tmr_registers(0)(590) and tmr_registers(1)(590)) or                                            
                            (tmr_registers(1)(590) and tmr_registers(2)(590)) or                                                       
                            (tmr_registers(0)(590) and tmr_registers(2)(590));                                                         
                                                                                                                                     
        global_tmr_voter(0)(591)  <=    (tmr_registers(0)(591) and tmr_registers(1)(591)) or                                            
                            (tmr_registers(1)(591) and tmr_registers(2)(591)) or                                                       
                            (tmr_registers(0)(591) and tmr_registers(2)(591));                                                         
                                                                                                                                     
        global_tmr_voter(0)(592)  <=    (tmr_registers(0)(592) and tmr_registers(1)(592)) or                                            
                            (tmr_registers(1)(592) and tmr_registers(2)(592)) or                                                       
                            (tmr_registers(0)(592) and tmr_registers(2)(592));                                                         
                                                                                                                                     
        global_tmr_voter(0)(593)  <=    (tmr_registers(0)(593) and tmr_registers(1)(593)) or                                            
                            (tmr_registers(1)(593) and tmr_registers(2)(593)) or                                                       
                            (tmr_registers(0)(593) and tmr_registers(2)(593));                                                         
                                                                                                                                     
        global_tmr_voter(0)(594)  <=    (tmr_registers(0)(594) and tmr_registers(1)(594)) or                                            
                            (tmr_registers(1)(594) and tmr_registers(2)(594)) or                                                       
                            (tmr_registers(0)(594) and tmr_registers(2)(594));                                                         
                                                                                                                                     
        global_tmr_voter(0)(595)  <=    (tmr_registers(0)(595) and tmr_registers(1)(595)) or                                            
                            (tmr_registers(1)(595) and tmr_registers(2)(595)) or                                                       
                            (tmr_registers(0)(595) and tmr_registers(2)(595));                                                         
                                                                                                                                     
        global_tmr_voter(0)(596)  <=    (tmr_registers(0)(596) and tmr_registers(1)(596)) or                                            
                            (tmr_registers(1)(596) and tmr_registers(2)(596)) or                                                       
                            (tmr_registers(0)(596) and tmr_registers(2)(596));                                                         
                                                                                                                                     
        global_tmr_voter(0)(597)  <=    (tmr_registers(0)(597) and tmr_registers(1)(597)) or                                            
                            (tmr_registers(1)(597) and tmr_registers(2)(597)) or                                                       
                            (tmr_registers(0)(597) and tmr_registers(2)(597));                                                         
                                                                                                                                     
        global_tmr_voter(0)(598)  <=    (tmr_registers(0)(598) and tmr_registers(1)(598)) or                                            
                            (tmr_registers(1)(598) and tmr_registers(2)(598)) or                                                       
                            (tmr_registers(0)(598) and tmr_registers(2)(598));                                                         
                                                                                                                                     
        global_tmr_voter(0)(599)  <=    (tmr_registers(0)(599) and tmr_registers(1)(599)) or                                            
                            (tmr_registers(1)(599) and tmr_registers(2)(599)) or                                                       
                            (tmr_registers(0)(599) and tmr_registers(2)(599));                                                         
                                                                                                                                     
        global_tmr_voter(0)(600)  <=    (tmr_registers(0)(600) and tmr_registers(1)(600)) or                                            
                            (tmr_registers(1)(600) and tmr_registers(2)(600)) or                                                       
                            (tmr_registers(0)(600) and tmr_registers(2)(600));                                                         
                                                                                                                                     
        global_tmr_voter(0)(601)  <=    (tmr_registers(0)(601) and tmr_registers(1)(601)) or                                            
                            (tmr_registers(1)(601) and tmr_registers(2)(601)) or                                                       
                            (tmr_registers(0)(601) and tmr_registers(2)(601));                                                         
                                                                                                                                     
        global_tmr_voter(0)(602)  <=    (tmr_registers(0)(602) and tmr_registers(1)(602)) or                                            
                            (tmr_registers(1)(602) and tmr_registers(2)(602)) or                                                       
                            (tmr_registers(0)(602) and tmr_registers(2)(602));                                                         
                                                                                                                                     
        global_tmr_voter(0)(603)  <=    (tmr_registers(0)(603) and tmr_registers(1)(603)) or                                            
                            (tmr_registers(1)(603) and tmr_registers(2)(603)) or                                                       
                            (tmr_registers(0)(603) and tmr_registers(2)(603));                                                         
                                                                                                                                     
        global_tmr_voter(0)(604)  <=    (tmr_registers(0)(604) and tmr_registers(1)(604)) or                                            
                            (tmr_registers(1)(604) and tmr_registers(2)(604)) or                                                       
                            (tmr_registers(0)(604) and tmr_registers(2)(604));                                                         
                                                                                                                                     
        global_tmr_voter(0)(605)  <=    (tmr_registers(0)(605) and tmr_registers(1)(605)) or                                            
                            (tmr_registers(1)(605) and tmr_registers(2)(605)) or                                                       
                            (tmr_registers(0)(605) and tmr_registers(2)(605));                                                         
                                                                                                                                     
        global_tmr_voter(0)(606)  <=    (tmr_registers(0)(606) and tmr_registers(1)(606)) or                                            
                            (tmr_registers(1)(606) and tmr_registers(2)(606)) or                                                       
                            (tmr_registers(0)(606) and tmr_registers(2)(606));                                                         
                                                                                                                                     
        global_tmr_voter(0)(607)  <=    (tmr_registers(0)(607) and tmr_registers(1)(607)) or                                            
                            (tmr_registers(1)(607) and tmr_registers(2)(607)) or                                                       
                            (tmr_registers(0)(607) and tmr_registers(2)(607));                                                         
                                                                                                                                     
        global_tmr_voter(0)(608)  <=    (tmr_registers(0)(608) and tmr_registers(1)(608)) or                                            
                            (tmr_registers(1)(608) and tmr_registers(2)(608)) or                                                       
                            (tmr_registers(0)(608) and tmr_registers(2)(608));                                                         
                                                                                                                                     
        global_tmr_voter(0)(609)  <=    (tmr_registers(0)(609) and tmr_registers(1)(609)) or                                            
                            (tmr_registers(1)(609) and tmr_registers(2)(609)) or                                                       
                            (tmr_registers(0)(609) and tmr_registers(2)(609));                                                         
                                                                                                                                     
        global_tmr_voter(0)(610)  <=    (tmr_registers(0)(610) and tmr_registers(1)(610)) or                                            
                            (tmr_registers(1)(610) and tmr_registers(2)(610)) or                                                       
                            (tmr_registers(0)(610) and tmr_registers(2)(610));                                                         
                                                                                                                                     
        global_tmr_voter(0)(611)  <=    (tmr_registers(0)(611) and tmr_registers(1)(611)) or                                            
                            (tmr_registers(1)(611) and tmr_registers(2)(611)) or                                                       
                            (tmr_registers(0)(611) and tmr_registers(2)(611));                                                         
                                                                                                                                     
        global_tmr_voter(0)(612)  <=    (tmr_registers(0)(612) and tmr_registers(1)(612)) or                                            
                            (tmr_registers(1)(612) and tmr_registers(2)(612)) or                                                       
                            (tmr_registers(0)(612) and tmr_registers(2)(612));                                                         
                                                                                                                                     
        global_tmr_voter(0)(613)  <=    (tmr_registers(0)(613) and tmr_registers(1)(613)) or                                            
                            (tmr_registers(1)(613) and tmr_registers(2)(613)) or                                                       
                            (tmr_registers(0)(613) and tmr_registers(2)(613));                                                         
                                                                                                                                     
        global_tmr_voter(0)(614)  <=    (tmr_registers(0)(614) and tmr_registers(1)(614)) or                                            
                            (tmr_registers(1)(614) and tmr_registers(2)(614)) or                                                       
                            (tmr_registers(0)(614) and tmr_registers(2)(614));                                                         
                                                                                                                                     
        global_tmr_voter(0)(615)  <=    (tmr_registers(0)(615) and tmr_registers(1)(615)) or                                            
                            (tmr_registers(1)(615) and tmr_registers(2)(615)) or                                                       
                            (tmr_registers(0)(615) and tmr_registers(2)(615));                                                         
                                                                                                                                     
        global_tmr_voter(0)(616)  <=    (tmr_registers(0)(616) and tmr_registers(1)(616)) or                                            
                            (tmr_registers(1)(616) and tmr_registers(2)(616)) or                                                       
                            (tmr_registers(0)(616) and tmr_registers(2)(616));                                                         
                                                                                                                                     
        global_tmr_voter(0)(617)  <=    (tmr_registers(0)(617) and tmr_registers(1)(617)) or                                            
                            (tmr_registers(1)(617) and tmr_registers(2)(617)) or                                                       
                            (tmr_registers(0)(617) and tmr_registers(2)(617));                                                         
                                                                                                                                     
        global_tmr_voter(0)(618)  <=    (tmr_registers(0)(618) and tmr_registers(1)(618)) or                                            
                            (tmr_registers(1)(618) and tmr_registers(2)(618)) or                                                       
                            (tmr_registers(0)(618) and tmr_registers(2)(618));                                                         
                                                                                                                                     
        global_tmr_voter(0)(619)  <=    (tmr_registers(0)(619) and tmr_registers(1)(619)) or                                            
                            (tmr_registers(1)(619) and tmr_registers(2)(619)) or                                                       
                            (tmr_registers(0)(619) and tmr_registers(2)(619));                                                         
                                                                                                                                     
        global_tmr_voter(0)(620)  <=    (tmr_registers(0)(620) and tmr_registers(1)(620)) or                                            
                            (tmr_registers(1)(620) and tmr_registers(2)(620)) or                                                       
                            (tmr_registers(0)(620) and tmr_registers(2)(620));                                                         
                                                                                                                                     
        global_tmr_voter(0)(621)  <=    (tmr_registers(0)(621) and tmr_registers(1)(621)) or                                            
                            (tmr_registers(1)(621) and tmr_registers(2)(621)) or                                                       
                            (tmr_registers(0)(621) and tmr_registers(2)(621));                                                         
                                                                                                                                     
        global_tmr_voter(0)(622)  <=    (tmr_registers(0)(622) and tmr_registers(1)(622)) or                                            
                            (tmr_registers(1)(622) and tmr_registers(2)(622)) or                                                       
                            (tmr_registers(0)(622) and tmr_registers(2)(622));                                                         
                                                                                                                                     
        global_tmr_voter(0)(623)  <=    (tmr_registers(0)(623) and tmr_registers(1)(623)) or                                            
                            (tmr_registers(1)(623) and tmr_registers(2)(623)) or                                                       
                            (tmr_registers(0)(623) and tmr_registers(2)(623));                                                         
                                                                                                                                     
        global_tmr_voter(0)(624)  <=    (tmr_registers(0)(624) and tmr_registers(1)(624)) or                                            
                            (tmr_registers(1)(624) and tmr_registers(2)(624)) or                                                       
                            (tmr_registers(0)(624) and tmr_registers(2)(624));                                                         
                                                                                                                                     
        global_tmr_voter(0)(625)  <=    (tmr_registers(0)(625) and tmr_registers(1)(625)) or                                            
                            (tmr_registers(1)(625) and tmr_registers(2)(625)) or                                                       
                            (tmr_registers(0)(625) and tmr_registers(2)(625));                                                         
                                                                                                                                     
        global_tmr_voter(0)(626)  <=    (tmr_registers(0)(626) and tmr_registers(1)(626)) or                                            
                            (tmr_registers(1)(626) and tmr_registers(2)(626)) or                                                       
                            (tmr_registers(0)(626) and tmr_registers(2)(626));                                                         
                                                                                                                                     
        global_tmr_voter(0)(627)  <=    (tmr_registers(0)(627) and tmr_registers(1)(627)) or                                            
                            (tmr_registers(1)(627) and tmr_registers(2)(627)) or                                                       
                            (tmr_registers(0)(627) and tmr_registers(2)(627));                                                         
                                                                                                                                     
        global_tmr_voter(0)(628)  <=    (tmr_registers(0)(628) and tmr_registers(1)(628)) or                                            
                            (tmr_registers(1)(628) and tmr_registers(2)(628)) or                                                       
                            (tmr_registers(0)(628) and tmr_registers(2)(628));                                                         
                                                                                                                                     
        global_tmr_voter(0)(629)  <=    (tmr_registers(0)(629) and tmr_registers(1)(629)) or                                            
                            (tmr_registers(1)(629) and tmr_registers(2)(629)) or                                                       
                            (tmr_registers(0)(629) and tmr_registers(2)(629));                                                         
                                                                                                                                     
        global_tmr_voter(0)(630)  <=    (tmr_registers(0)(630) and tmr_registers(1)(630)) or                                            
                            (tmr_registers(1)(630) and tmr_registers(2)(630)) or                                                       
                            (tmr_registers(0)(630) and tmr_registers(2)(630));                                                         
                                                                                                                                     
        global_tmr_voter(0)(631)  <=    (tmr_registers(0)(631) and tmr_registers(1)(631)) or                                            
                            (tmr_registers(1)(631) and tmr_registers(2)(631)) or                                                       
                            (tmr_registers(0)(631) and tmr_registers(2)(631));                                                         
                                                                                                                                     
        global_tmr_voter(0)(632)  <=    (tmr_registers(0)(632) and tmr_registers(1)(632)) or                                            
                            (tmr_registers(1)(632) and tmr_registers(2)(632)) or                                                       
                            (tmr_registers(0)(632) and tmr_registers(2)(632));                                                         
                                                                                                                                     
        global_tmr_voter(0)(633)  <=    (tmr_registers(0)(633) and tmr_registers(1)(633)) or                                            
                            (tmr_registers(1)(633) and tmr_registers(2)(633)) or                                                       
                            (tmr_registers(0)(633) and tmr_registers(2)(633));                                                         
                                                                                                                                     
        global_tmr_voter(0)(634)  <=    (tmr_registers(0)(634) and tmr_registers(1)(634)) or                                            
                            (tmr_registers(1)(634) and tmr_registers(2)(634)) or                                                       
                            (tmr_registers(0)(634) and tmr_registers(2)(634));                                                         
                                                                                                                                     
        global_tmr_voter(0)(635)  <=    (tmr_registers(0)(635) and tmr_registers(1)(635)) or                                            
                            (tmr_registers(1)(635) and tmr_registers(2)(635)) or                                                       
                            (tmr_registers(0)(635) and tmr_registers(2)(635));                                                         
                                                                                                                                     
        global_tmr_voter(0)(636)  <=    (tmr_registers(0)(636) and tmr_registers(1)(636)) or                                            
                            (tmr_registers(1)(636) and tmr_registers(2)(636)) or                                                       
                            (tmr_registers(0)(636) and tmr_registers(2)(636));                                                         
                                                                                                                                     
        global_tmr_voter(0)(637)  <=    (tmr_registers(0)(637) and tmr_registers(1)(637)) or                                            
                            (tmr_registers(1)(637) and tmr_registers(2)(637)) or                                                       
                            (tmr_registers(0)(637) and tmr_registers(2)(637));                                                         
                                                                                                                                     
        global_tmr_voter(0)(638)  <=    (tmr_registers(0)(638) and tmr_registers(1)(638)) or                                            
                            (tmr_registers(1)(638) and tmr_registers(2)(638)) or                                                       
                            (tmr_registers(0)(638) and tmr_registers(2)(638));                                                         
                                                                                                                                     
        global_tmr_voter(0)(639)  <=    (tmr_registers(0)(639) and tmr_registers(1)(639)) or                                            
                            (tmr_registers(1)(639) and tmr_registers(2)(639)) or                                                       
                            (tmr_registers(0)(639) and tmr_registers(2)(639));                                                         
                                                                                                                                     
        global_tmr_voter(0)(640)  <=    (tmr_registers(0)(640) and tmr_registers(1)(640)) or                                            
                            (tmr_registers(1)(640) and tmr_registers(2)(640)) or                                                       
                            (tmr_registers(0)(640) and tmr_registers(2)(640));                                                         
                                                                                                                                     
        global_tmr_voter(0)(641)  <=    (tmr_registers(0)(641) and tmr_registers(1)(641)) or                                            
                            (tmr_registers(1)(641) and tmr_registers(2)(641)) or                                                       
                            (tmr_registers(0)(641) and tmr_registers(2)(641));                                                         
                                                                                                                                     
        global_tmr_voter(0)(642)  <=    (tmr_registers(0)(642) and tmr_registers(1)(642)) or                                            
                            (tmr_registers(1)(642) and tmr_registers(2)(642)) or                                                       
                            (tmr_registers(0)(642) and tmr_registers(2)(642));                                                         
                                                                                                                                     
        global_tmr_voter(0)(643)  <=    (tmr_registers(0)(643) and tmr_registers(1)(643)) or                                            
                            (tmr_registers(1)(643) and tmr_registers(2)(643)) or                                                       
                            (tmr_registers(0)(643) and tmr_registers(2)(643));                                                         
                                                                                                                                     
        global_tmr_voter(0)(644)  <=    (tmr_registers(0)(644) and tmr_registers(1)(644)) or                                            
                            (tmr_registers(1)(644) and tmr_registers(2)(644)) or                                                       
                            (tmr_registers(0)(644) and tmr_registers(2)(644));                                                         
                                                                                                                                     
        global_tmr_voter(0)(645)  <=    (tmr_registers(0)(645) and tmr_registers(1)(645)) or                                            
                            (tmr_registers(1)(645) and tmr_registers(2)(645)) or                                                       
                            (tmr_registers(0)(645) and tmr_registers(2)(645));                                                         
                                                                                                                                     
        global_tmr_voter(0)(646)  <=    (tmr_registers(0)(646) and tmr_registers(1)(646)) or                                            
                            (tmr_registers(1)(646) and tmr_registers(2)(646)) or                                                       
                            (tmr_registers(0)(646) and tmr_registers(2)(646));                                                         
                                                                                                                                     
        global_tmr_voter(0)(647)  <=    (tmr_registers(0)(647) and tmr_registers(1)(647)) or                                            
                            (tmr_registers(1)(647) and tmr_registers(2)(647)) or                                                       
                            (tmr_registers(0)(647) and tmr_registers(2)(647));                                                         
                                                                                                                                     
        global_tmr_voter(0)(648)  <=    (tmr_registers(0)(648) and tmr_registers(1)(648)) or                                            
                            (tmr_registers(1)(648) and tmr_registers(2)(648)) or                                                       
                            (tmr_registers(0)(648) and tmr_registers(2)(648));                                                         
                                                                                                                                     
        global_tmr_voter(0)(649)  <=    (tmr_registers(0)(649) and tmr_registers(1)(649)) or                                            
                            (tmr_registers(1)(649) and tmr_registers(2)(649)) or                                                       
                            (tmr_registers(0)(649) and tmr_registers(2)(649));                                                         
                                                                                                                                     
        global_tmr_voter(0)(650)  <=    (tmr_registers(0)(650) and tmr_registers(1)(650)) or                                            
                            (tmr_registers(1)(650) and tmr_registers(2)(650)) or                                                       
                            (tmr_registers(0)(650) and tmr_registers(2)(650));                                                         
                                                                                                                                     
        global_tmr_voter(0)(651)  <=    (tmr_registers(0)(651) and tmr_registers(1)(651)) or                                            
                            (tmr_registers(1)(651) and tmr_registers(2)(651)) or                                                       
                            (tmr_registers(0)(651) and tmr_registers(2)(651));                                                         
                                                                                                                                     
        global_tmr_voter(0)(652)  <=    (tmr_registers(0)(652) and tmr_registers(1)(652)) or                                            
                            (tmr_registers(1)(652) and tmr_registers(2)(652)) or                                                       
                            (tmr_registers(0)(652) and tmr_registers(2)(652));                                                         
                                                                                                                                     
        global_tmr_voter(0)(653)  <=    (tmr_registers(0)(653) and tmr_registers(1)(653)) or                                            
                            (tmr_registers(1)(653) and tmr_registers(2)(653)) or                                                       
                            (tmr_registers(0)(653) and tmr_registers(2)(653));                                                         
                                                                                                                                     
        global_tmr_voter(0)(654)  <=    (tmr_registers(0)(654) and tmr_registers(1)(654)) or                                            
                            (tmr_registers(1)(654) and tmr_registers(2)(654)) or                                                       
                            (tmr_registers(0)(654) and tmr_registers(2)(654));                                                         
                                                                                                                                     
        global_tmr_voter(0)(655)  <=    (tmr_registers(0)(655) and tmr_registers(1)(655)) or                                            
                            (tmr_registers(1)(655) and tmr_registers(2)(655)) or                                                       
                            (tmr_registers(0)(655) and tmr_registers(2)(655));                                                         
                                                                                                                                     
        global_tmr_voter(0)(656)  <=    (tmr_registers(0)(656) and tmr_registers(1)(656)) or                                            
                            (tmr_registers(1)(656) and tmr_registers(2)(656)) or                                                       
                            (tmr_registers(0)(656) and tmr_registers(2)(656));                                                         
                                                                                                                                     
        global_tmr_voter(0)(657)  <=    (tmr_registers(0)(657) and tmr_registers(1)(657)) or                                            
                            (tmr_registers(1)(657) and tmr_registers(2)(657)) or                                                       
                            (tmr_registers(0)(657) and tmr_registers(2)(657));                                                         
                                                                                                                                     
        global_tmr_voter(0)(658)  <=    (tmr_registers(0)(658) and tmr_registers(1)(658)) or                                            
                            (tmr_registers(1)(658) and tmr_registers(2)(658)) or                                                       
                            (tmr_registers(0)(658) and tmr_registers(2)(658));                                                         
                                                                                                                                     
        global_tmr_voter(0)(659)  <=    (tmr_registers(0)(659) and tmr_registers(1)(659)) or                                            
                            (tmr_registers(1)(659) and tmr_registers(2)(659)) or                                                       
                            (tmr_registers(0)(659) and tmr_registers(2)(659));                                                         
                                                                                                                                     
        global_tmr_voter(0)(660)  <=    (tmr_registers(0)(660) and tmr_registers(1)(660)) or                                            
                            (tmr_registers(1)(660) and tmr_registers(2)(660)) or                                                       
                            (tmr_registers(0)(660) and tmr_registers(2)(660));                                                         
                                                                                                                                     
        global_tmr_voter(0)(661)  <=    (tmr_registers(0)(661) and tmr_registers(1)(661)) or                                            
                            (tmr_registers(1)(661) and tmr_registers(2)(661)) or                                                       
                            (tmr_registers(0)(661) and tmr_registers(2)(661));                                                         
                                                                                                                                     
        global_tmr_voter(0)(662)  <=    (tmr_registers(0)(662) and tmr_registers(1)(662)) or                                            
                            (tmr_registers(1)(662) and tmr_registers(2)(662)) or                                                       
                            (tmr_registers(0)(662) and tmr_registers(2)(662));                                                         
                                                                                                                                     
        global_tmr_voter(0)(663)  <=    (tmr_registers(0)(663) and tmr_registers(1)(663)) or                                            
                            (tmr_registers(1)(663) and tmr_registers(2)(663)) or                                                       
                            (tmr_registers(0)(663) and tmr_registers(2)(663));                                                         
                                                                                                                                     
        global_tmr_voter(0)(664)  <=    (tmr_registers(0)(664) and tmr_registers(1)(664)) or                                            
                            (tmr_registers(1)(664) and tmr_registers(2)(664)) or                                                       
                            (tmr_registers(0)(664) and tmr_registers(2)(664));                                                         
                                                                                                                                     
        global_tmr_voter(0)(665)  <=    (tmr_registers(0)(665) and tmr_registers(1)(665)) or                                            
                            (tmr_registers(1)(665) and tmr_registers(2)(665)) or                                                       
                            (tmr_registers(0)(665) and tmr_registers(2)(665));                                                         
                                                                                                                                     
        global_tmr_voter(0)(666)  <=    (tmr_registers(0)(666) and tmr_registers(1)(666)) or                                            
                            (tmr_registers(1)(666) and tmr_registers(2)(666)) or                                                       
                            (tmr_registers(0)(666) and tmr_registers(2)(666));                                                         
                                                                                                                                     
        global_tmr_voter(0)(667)  <=    (tmr_registers(0)(667) and tmr_registers(1)(667)) or                                            
                            (tmr_registers(1)(667) and tmr_registers(2)(667)) or                                                       
                            (tmr_registers(0)(667) and tmr_registers(2)(667));                                                         
                                                                                                                                     
        global_tmr_voter(0)(668)  <=    (tmr_registers(0)(668) and tmr_registers(1)(668)) or                                            
                            (tmr_registers(1)(668) and tmr_registers(2)(668)) or                                                       
                            (tmr_registers(0)(668) and tmr_registers(2)(668));                                                         
                                                                                                                                     
        global_tmr_voter(0)(669)  <=    (tmr_registers(0)(669) and tmr_registers(1)(669)) or                                            
                            (tmr_registers(1)(669) and tmr_registers(2)(669)) or                                                       
                            (tmr_registers(0)(669) and tmr_registers(2)(669));                                                         
                                                                                                                                     
        global_tmr_voter(0)(670)  <=    (tmr_registers(0)(670) and tmr_registers(1)(670)) or                                            
                            (tmr_registers(1)(670) and tmr_registers(2)(670)) or                                                       
                            (tmr_registers(0)(670) and tmr_registers(2)(670));                                                         
                                                                                                                                     
        global_tmr_voter(0)(671)  <=    (tmr_registers(0)(671) and tmr_registers(1)(671)) or                                            
                            (tmr_registers(1)(671) and tmr_registers(2)(671)) or                                                       
                            (tmr_registers(0)(671) and tmr_registers(2)(671));                                                         
                                                                                                                                     
        global_tmr_voter(0)(672)  <=    (tmr_registers(0)(672) and tmr_registers(1)(672)) or                                            
                            (tmr_registers(1)(672) and tmr_registers(2)(672)) or                                                       
                            (tmr_registers(0)(672) and tmr_registers(2)(672));                                                         
                                                                                                                                     
        global_tmr_voter(0)(673)  <=    (tmr_registers(0)(673) and tmr_registers(1)(673)) or                                            
                            (tmr_registers(1)(673) and tmr_registers(2)(673)) or                                                       
                            (tmr_registers(0)(673) and tmr_registers(2)(673));                                                         
                                                                                                                                     
        global_tmr_voter(0)(674)  <=    (tmr_registers(0)(674) and tmr_registers(1)(674)) or                                            
                            (tmr_registers(1)(674) and tmr_registers(2)(674)) or                                                       
                            (tmr_registers(0)(674) and tmr_registers(2)(674));                                                         
                                                                                                                                     
        global_tmr_voter(0)(675)  <=    (tmr_registers(0)(675) and tmr_registers(1)(675)) or                                            
                            (tmr_registers(1)(675) and tmr_registers(2)(675)) or                                                       
                            (tmr_registers(0)(675) and tmr_registers(2)(675));                                                         
                                                                                                                                     
        global_tmr_voter(0)(676)  <=    (tmr_registers(0)(676) and tmr_registers(1)(676)) or                                            
                            (tmr_registers(1)(676) and tmr_registers(2)(676)) or                                                       
                            (tmr_registers(0)(676) and tmr_registers(2)(676));                                                         
                                                                                                                                     
        global_tmr_voter(0)(677)  <=    (tmr_registers(0)(677) and tmr_registers(1)(677)) or                                            
                            (tmr_registers(1)(677) and tmr_registers(2)(677)) or                                                       
                            (tmr_registers(0)(677) and tmr_registers(2)(677));                                                         
                                                                                                                                     
        global_tmr_voter(0)(678)  <=    (tmr_registers(0)(678) and tmr_registers(1)(678)) or                                            
                            (tmr_registers(1)(678) and tmr_registers(2)(678)) or                                                       
                            (tmr_registers(0)(678) and tmr_registers(2)(678));                                                         
                                                                                                                                     
        global_tmr_voter(0)(679)  <=    (tmr_registers(0)(679) and tmr_registers(1)(679)) or                                            
                            (tmr_registers(1)(679) and tmr_registers(2)(679)) or                                                       
                            (tmr_registers(0)(679) and tmr_registers(2)(679));                                                         
                                                                                                                                     
        global_tmr_voter(0)(680)  <=    (tmr_registers(0)(680) and tmr_registers(1)(680)) or                                            
                            (tmr_registers(1)(680) and tmr_registers(2)(680)) or                                                       
                            (tmr_registers(0)(680) and tmr_registers(2)(680));                                                         
                                                                                                                                     
        global_tmr_voter(0)(681)  <=    (tmr_registers(0)(681) and tmr_registers(1)(681)) or                                            
                            (tmr_registers(1)(681) and tmr_registers(2)(681)) or                                                       
                            (tmr_registers(0)(681) and tmr_registers(2)(681));                                                         
                                                                                                                                     
        global_tmr_voter(0)(682)  <=    (tmr_registers(0)(682) and tmr_registers(1)(682)) or                                            
                            (tmr_registers(1)(682) and tmr_registers(2)(682)) or                                                       
                            (tmr_registers(0)(682) and tmr_registers(2)(682));                                                         
                                                                                                                                     
        global_tmr_voter(0)(683)  <=    (tmr_registers(0)(683) and tmr_registers(1)(683)) or                                            
                            (tmr_registers(1)(683) and tmr_registers(2)(683)) or                                                       
                            (tmr_registers(0)(683) and tmr_registers(2)(683));                                                         
                                                                                                                                     
        global_tmr_voter(0)(684)  <=    (tmr_registers(0)(684) and tmr_registers(1)(684)) or                                            
                            (tmr_registers(1)(684) and tmr_registers(2)(684)) or                                                       
                            (tmr_registers(0)(684) and tmr_registers(2)(684));                                                         
                                                                                                                                     
        global_tmr_voter(0)(685)  <=    (tmr_registers(0)(685) and tmr_registers(1)(685)) or                                            
                            (tmr_registers(1)(685) and tmr_registers(2)(685)) or                                                       
                            (tmr_registers(0)(685) and tmr_registers(2)(685));                                                         
                                                                                                                                     
        global_tmr_voter(0)(686)  <=    (tmr_registers(0)(686) and tmr_registers(1)(686)) or                                            
                            (tmr_registers(1)(686) and tmr_registers(2)(686)) or                                                       
                            (tmr_registers(0)(686) and tmr_registers(2)(686));                                                         
                                                                                                                                     
        global_tmr_voter(0)(687)  <=    (tmr_registers(0)(687) and tmr_registers(1)(687)) or                                            
                            (tmr_registers(1)(687) and tmr_registers(2)(687)) or                                                       
                            (tmr_registers(0)(687) and tmr_registers(2)(687));                                                         
                                                                                                                                     
        global_tmr_voter(0)(688)  <=    (tmr_registers(0)(688) and tmr_registers(1)(688)) or                                            
                            (tmr_registers(1)(688) and tmr_registers(2)(688)) or                                                       
                            (tmr_registers(0)(688) and tmr_registers(2)(688));                                                         
                                                                                                                                     
        global_tmr_voter(0)(689)  <=    (tmr_registers(0)(689) and tmr_registers(1)(689)) or                                            
                            (tmr_registers(1)(689) and tmr_registers(2)(689)) or                                                       
                            (tmr_registers(0)(689) and tmr_registers(2)(689));                                                         
                                                                                                                                     
        global_tmr_voter(0)(690)  <=    (tmr_registers(0)(690) and tmr_registers(1)(690)) or                                            
                            (tmr_registers(1)(690) and tmr_registers(2)(690)) or                                                       
                            (tmr_registers(0)(690) and tmr_registers(2)(690));                                                         
                                                                                                                                     
        global_tmr_voter(0)(691)  <=    (tmr_registers(0)(691) and tmr_registers(1)(691)) or                                            
                            (tmr_registers(1)(691) and tmr_registers(2)(691)) or                                                       
                            (tmr_registers(0)(691) and tmr_registers(2)(691));                                                         
                                                                                                                                     
        global_tmr_voter(0)(692)  <=    (tmr_registers(0)(692) and tmr_registers(1)(692)) or                                            
                            (tmr_registers(1)(692) and tmr_registers(2)(692)) or                                                       
                            (tmr_registers(0)(692) and tmr_registers(2)(692));                                                         
                                                                                                                                     
        global_tmr_voter(0)(693)  <=    (tmr_registers(0)(693) and tmr_registers(1)(693)) or                                            
                            (tmr_registers(1)(693) and tmr_registers(2)(693)) or                                                       
                            (tmr_registers(0)(693) and tmr_registers(2)(693));                                                         
                                                                                                                                     
        global_tmr_voter(0)(694)  <=    (tmr_registers(0)(694) and tmr_registers(1)(694)) or                                            
                            (tmr_registers(1)(694) and tmr_registers(2)(694)) or                                                       
                            (tmr_registers(0)(694) and tmr_registers(2)(694));                                                         
                                                                                                                                     
        global_tmr_voter(0)(695)  <=    (tmr_registers(0)(695) and tmr_registers(1)(695)) or                                            
                            (tmr_registers(1)(695) and tmr_registers(2)(695)) or                                                       
                            (tmr_registers(0)(695) and tmr_registers(2)(695));                                                         
                                                                                                                                     
        global_tmr_voter(0)(696)  <=    (tmr_registers(0)(696) and tmr_registers(1)(696)) or                                            
                            (tmr_registers(1)(696) and tmr_registers(2)(696)) or                                                       
                            (tmr_registers(0)(696) and tmr_registers(2)(696));                                                         
                                                                                                                                     
        global_tmr_voter(0)(697)  <=    (tmr_registers(0)(697) and tmr_registers(1)(697)) or                                            
                            (tmr_registers(1)(697) and tmr_registers(2)(697)) or                                                       
                            (tmr_registers(0)(697) and tmr_registers(2)(697));                                                         
                                                                                                                                     
        global_tmr_voter(0)(698)  <=    (tmr_registers(0)(698) and tmr_registers(1)(698)) or                                            
                            (tmr_registers(1)(698) and tmr_registers(2)(698)) or                                                       
                            (tmr_registers(0)(698) and tmr_registers(2)(698));                                                         
                                                                                                                                     
        global_tmr_voter(0)(699)  <=    (tmr_registers(0)(699) and tmr_registers(1)(699)) or                                            
                            (tmr_registers(1)(699) and tmr_registers(2)(699)) or                                                       
                            (tmr_registers(0)(699) and tmr_registers(2)(699));                                                         
                                                                                                                                     
        global_tmr_voter(0)(700)  <=    (tmr_registers(0)(700) and tmr_registers(1)(700)) or                                            
                            (tmr_registers(1)(700) and tmr_registers(2)(700)) or                                                       
                            (tmr_registers(0)(700) and tmr_registers(2)(700));                                                         
                                                                                                                                     
        global_tmr_voter(0)(701)  <=    (tmr_registers(0)(701) and tmr_registers(1)(701)) or                                            
                            (tmr_registers(1)(701) and tmr_registers(2)(701)) or                                                       
                            (tmr_registers(0)(701) and tmr_registers(2)(701));                                                         
                                                                                                                                     
        global_tmr_voter(0)(702)  <=    (tmr_registers(0)(702) and tmr_registers(1)(702)) or                                            
                            (tmr_registers(1)(702) and tmr_registers(2)(702)) or                                                       
                            (tmr_registers(0)(702) and tmr_registers(2)(702));                                                         
                                                                                                                                     
        global_tmr_voter(0)(703)  <=    (tmr_registers(0)(703) and tmr_registers(1)(703)) or                                            
                            (tmr_registers(1)(703) and tmr_registers(2)(703)) or                                                       
                            (tmr_registers(0)(703) and tmr_registers(2)(703));                                                         
                                                                                                                                     
        global_tmr_voter(0)(704)  <=    (tmr_registers(0)(704) and tmr_registers(1)(704)) or                                            
                            (tmr_registers(1)(704) and tmr_registers(2)(704)) or                                                       
                            (tmr_registers(0)(704) and tmr_registers(2)(704));                                                         
                                                                                                                                     
        global_tmr_voter(0)(705)  <=    (tmr_registers(0)(705) and tmr_registers(1)(705)) or                                            
                            (tmr_registers(1)(705) and tmr_registers(2)(705)) or                                                       
                            (tmr_registers(0)(705) and tmr_registers(2)(705));                                                         
                                                                                                                                     
        global_tmr_voter(0)(706)  <=    (tmr_registers(0)(706) and tmr_registers(1)(706)) or                                            
                            (tmr_registers(1)(706) and tmr_registers(2)(706)) or                                                       
                            (tmr_registers(0)(706) and tmr_registers(2)(706));                                                         
                                                                                                                                     
        global_tmr_voter(0)(707)  <=    (tmr_registers(0)(707) and tmr_registers(1)(707)) or                                            
                            (tmr_registers(1)(707) and tmr_registers(2)(707)) or                                                       
                            (tmr_registers(0)(707) and tmr_registers(2)(707));                                                         
                                                                                                                                     
        global_tmr_voter(0)(708)  <=    (tmr_registers(0)(708) and tmr_registers(1)(708)) or                                            
                            (tmr_registers(1)(708) and tmr_registers(2)(708)) or                                                       
                            (tmr_registers(0)(708) and tmr_registers(2)(708));                                                         
                                                                                                                                     
        global_tmr_voter(0)(709)  <=    (tmr_registers(0)(709) and tmr_registers(1)(709)) or                                            
                            (tmr_registers(1)(709) and tmr_registers(2)(709)) or                                                       
                            (tmr_registers(0)(709) and tmr_registers(2)(709));                                                         
                                                                                                                                     
        global_tmr_voter(0)(710)  <=    (tmr_registers(0)(710) and tmr_registers(1)(710)) or                                            
                            (tmr_registers(1)(710) and tmr_registers(2)(710)) or                                                       
                            (tmr_registers(0)(710) and tmr_registers(2)(710));                                                         
                                                                                                                                     
        global_tmr_voter(0)(711)  <=    (tmr_registers(0)(711) and tmr_registers(1)(711)) or                                            
                            (tmr_registers(1)(711) and tmr_registers(2)(711)) or                                                       
                            (tmr_registers(0)(711) and tmr_registers(2)(711));                                                         
                                                                                                                                     
        global_tmr_voter(0)(712)  <=    (tmr_registers(0)(712) and tmr_registers(1)(712)) or                                            
                            (tmr_registers(1)(712) and tmr_registers(2)(712)) or                                                       
                            (tmr_registers(0)(712) and tmr_registers(2)(712));                                                         
                                                                                                                                     
        global_tmr_voter(0)(713)  <=    (tmr_registers(0)(713) and tmr_registers(1)(713)) or                                            
                            (tmr_registers(1)(713) and tmr_registers(2)(713)) or                                                       
                            (tmr_registers(0)(713) and tmr_registers(2)(713));                                                         
                                                                                                                                     
        global_tmr_voter(0)(714)  <=    (tmr_registers(0)(714) and tmr_registers(1)(714)) or                                            
                            (tmr_registers(1)(714) and tmr_registers(2)(714)) or                                                       
                            (tmr_registers(0)(714) and tmr_registers(2)(714));                                                         
                                                                                                                                     
        global_tmr_voter(0)(715)  <=    (tmr_registers(0)(715) and tmr_registers(1)(715)) or                                            
                            (tmr_registers(1)(715) and tmr_registers(2)(715)) or                                                       
                            (tmr_registers(0)(715) and tmr_registers(2)(715));                                                         
                                                                                                                                     
        global_tmr_voter(0)(716)  <=    (tmr_registers(0)(716) and tmr_registers(1)(716)) or                                            
                            (tmr_registers(1)(716) and tmr_registers(2)(716)) or                                                       
                            (tmr_registers(0)(716) and tmr_registers(2)(716));                                                         
                                                                                                                                     
        global_tmr_voter(0)(717)  <=    (tmr_registers(0)(717) and tmr_registers(1)(717)) or                                            
                            (tmr_registers(1)(717) and tmr_registers(2)(717)) or                                                       
                            (tmr_registers(0)(717) and tmr_registers(2)(717));                                                         
                                                                                                                                     
        global_tmr_voter(0)(718)  <=    (tmr_registers(0)(718) and tmr_registers(1)(718)) or                                            
                            (tmr_registers(1)(718) and tmr_registers(2)(718)) or                                                       
                            (tmr_registers(0)(718) and tmr_registers(2)(718));                                                         
                                                                                                                                     
        global_tmr_voter(0)(719)  <=    (tmr_registers(0)(719) and tmr_registers(1)(719)) or                                            
                            (tmr_registers(1)(719) and tmr_registers(2)(719)) or                                                       
                            (tmr_registers(0)(719) and tmr_registers(2)(719));                                                         
                                                                                                                                     
        global_tmr_voter(0)(720)  <=    (tmr_registers(0)(720) and tmr_registers(1)(720)) or                                            
                            (tmr_registers(1)(720) and tmr_registers(2)(720)) or                                                       
                            (tmr_registers(0)(720) and tmr_registers(2)(720));                                                         
                                                                                                                                     
        global_tmr_voter(0)(721)  <=    (tmr_registers(0)(721) and tmr_registers(1)(721)) or                                            
                            (tmr_registers(1)(721) and tmr_registers(2)(721)) or                                                       
                            (tmr_registers(0)(721) and tmr_registers(2)(721));                                                         
                                                                                                                                     
        global_tmr_voter(0)(722)  <=    (tmr_registers(0)(722) and tmr_registers(1)(722)) or                                            
                            (tmr_registers(1)(722) and tmr_registers(2)(722)) or                                                       
                            (tmr_registers(0)(722) and tmr_registers(2)(722));                                                         
                                                                                                                                     
        global_tmr_voter(0)(723)  <=    (tmr_registers(0)(723) and tmr_registers(1)(723)) or                                            
                            (tmr_registers(1)(723) and tmr_registers(2)(723)) or                                                       
                            (tmr_registers(0)(723) and tmr_registers(2)(723));                                                         
                                                                                                                                     
        global_tmr_voter(0)(724)  <=    (tmr_registers(0)(724) and tmr_registers(1)(724)) or                                            
                            (tmr_registers(1)(724) and tmr_registers(2)(724)) or                                                       
                            (tmr_registers(0)(724) and tmr_registers(2)(724));                                                         
                                                                                                                                     
        global_tmr_voter(0)(725)  <=    (tmr_registers(0)(725) and tmr_registers(1)(725)) or                                            
                            (tmr_registers(1)(725) and tmr_registers(2)(725)) or                                                       
                            (tmr_registers(0)(725) and tmr_registers(2)(725));                                                         
                                                                                                                                     
        global_tmr_voter(0)(726)  <=    (tmr_registers(0)(726) and tmr_registers(1)(726)) or                                            
                            (tmr_registers(1)(726) and tmr_registers(2)(726)) or                                                       
                            (tmr_registers(0)(726) and tmr_registers(2)(726));                                                         
                                                                                                                                     
        global_tmr_voter(0)(727)  <=    (tmr_registers(0)(727) and tmr_registers(1)(727)) or                                            
                            (tmr_registers(1)(727) and tmr_registers(2)(727)) or                                                       
                            (tmr_registers(0)(727) and tmr_registers(2)(727));                                                         
                                                                                                                                     
        global_tmr_voter(0)(728)  <=    (tmr_registers(0)(728) and tmr_registers(1)(728)) or                                            
                            (tmr_registers(1)(728) and tmr_registers(2)(728)) or                                                       
                            (tmr_registers(0)(728) and tmr_registers(2)(728));                                                         
                                                                                                                                     
        global_tmr_voter(0)(729)  <=    (tmr_registers(0)(729) and tmr_registers(1)(729)) or                                            
                            (tmr_registers(1)(729) and tmr_registers(2)(729)) or                                                       
                            (tmr_registers(0)(729) and tmr_registers(2)(729));                                                         
                                                                                                                                     
        global_tmr_voter(0)(730)  <=    (tmr_registers(0)(730) and tmr_registers(1)(730)) or                                            
                            (tmr_registers(1)(730) and tmr_registers(2)(730)) or                                                       
                            (tmr_registers(0)(730) and tmr_registers(2)(730));                                                         
                                                                                                                                     
        global_tmr_voter(0)(731)  <=    (tmr_registers(0)(731) and tmr_registers(1)(731)) or                                            
                            (tmr_registers(1)(731) and tmr_registers(2)(731)) or                                                       
                            (tmr_registers(0)(731) and tmr_registers(2)(731));                                                         
                                                                                                                                     
        global_tmr_voter(0)(732)  <=    (tmr_registers(0)(732) and tmr_registers(1)(732)) or                                            
                            (tmr_registers(1)(732) and tmr_registers(2)(732)) or                                                       
                            (tmr_registers(0)(732) and tmr_registers(2)(732));                                                         
                                                                                                                                     
        global_tmr_voter(0)(733)  <=    (tmr_registers(0)(733) and tmr_registers(1)(733)) or                                            
                            (tmr_registers(1)(733) and tmr_registers(2)(733)) or                                                       
                            (tmr_registers(0)(733) and tmr_registers(2)(733));                                                         
                                                                                                                                     
        global_tmr_voter(0)(734)  <=    (tmr_registers(0)(734) and tmr_registers(1)(734)) or                                            
                            (tmr_registers(1)(734) and tmr_registers(2)(734)) or                                                       
                            (tmr_registers(0)(734) and tmr_registers(2)(734));                                                         
                                                                                                                                     
        global_tmr_voter(0)(735)  <=    (tmr_registers(0)(735) and tmr_registers(1)(735)) or                                            
                            (tmr_registers(1)(735) and tmr_registers(2)(735)) or                                                       
                            (tmr_registers(0)(735) and tmr_registers(2)(735));                                                         
                                                                                                                                     
        global_tmr_voter(0)(736)  <=    (tmr_registers(0)(736) and tmr_registers(1)(736)) or                                            
                            (tmr_registers(1)(736) and tmr_registers(2)(736)) or                                                       
                            (tmr_registers(0)(736) and tmr_registers(2)(736));                                                         
                                                                                                                                     
        global_tmr_voter(0)(737)  <=    (tmr_registers(0)(737) and tmr_registers(1)(737)) or                                            
                            (tmr_registers(1)(737) and tmr_registers(2)(737)) or                                                       
                            (tmr_registers(0)(737) and tmr_registers(2)(737));                                                         
                                                                                                                                     
        global_tmr_voter(0)(738)  <=    (tmr_registers(0)(738) and tmr_registers(1)(738)) or                                            
                            (tmr_registers(1)(738) and tmr_registers(2)(738)) or                                                       
                            (tmr_registers(0)(738) and tmr_registers(2)(738));                                                         
                                                                                                                                     
        global_tmr_voter(0)(739)  <=    (tmr_registers(0)(739) and tmr_registers(1)(739)) or                                            
                            (tmr_registers(1)(739) and tmr_registers(2)(739)) or                                                       
                            (tmr_registers(0)(739) and tmr_registers(2)(739));                                                         
                                                                                                                                     
        global_tmr_voter(0)(740)  <=    (tmr_registers(0)(740) and tmr_registers(1)(740)) or                                            
                            (tmr_registers(1)(740) and tmr_registers(2)(740)) or                                                       
                            (tmr_registers(0)(740) and tmr_registers(2)(740));                                                         
                                                                                                                                     
        global_tmr_voter(0)(741)  <=    (tmr_registers(0)(741) and tmr_registers(1)(741)) or                                            
                            (tmr_registers(1)(741) and tmr_registers(2)(741)) or                                                       
                            (tmr_registers(0)(741) and tmr_registers(2)(741));                                                         
                                                                                                                                     
        global_tmr_voter(0)(742)  <=    (tmr_registers(0)(742) and tmr_registers(1)(742)) or                                            
                            (tmr_registers(1)(742) and tmr_registers(2)(742)) or                                                       
                            (tmr_registers(0)(742) and tmr_registers(2)(742));                                                         
                                                                                                                                     
        global_tmr_voter(0)(743)  <=    (tmr_registers(0)(743) and tmr_registers(1)(743)) or                                            
                            (tmr_registers(1)(743) and tmr_registers(2)(743)) or                                                       
                            (tmr_registers(0)(743) and tmr_registers(2)(743));                                                         
                                                                                                                                     
        global_tmr_voter(0)(744)  <=    (tmr_registers(0)(744) and tmr_registers(1)(744)) or                                            
                            (tmr_registers(1)(744) and tmr_registers(2)(744)) or                                                       
                            (tmr_registers(0)(744) and tmr_registers(2)(744));                                                         
                                                                                                                                     
        global_tmr_voter(0)(745)  <=    (tmr_registers(0)(745) and tmr_registers(1)(745)) or                                            
                            (tmr_registers(1)(745) and tmr_registers(2)(745)) or                                                       
                            (tmr_registers(0)(745) and tmr_registers(2)(745));                                                         
                                                                                                                                     
        global_tmr_voter(0)(746)  <=    (tmr_registers(0)(746) and tmr_registers(1)(746)) or                                            
                            (tmr_registers(1)(746) and tmr_registers(2)(746)) or                                                       
                            (tmr_registers(0)(746) and tmr_registers(2)(746));                                                         
                                                                                                                                     
        global_tmr_voter(0)(747)  <=    (tmr_registers(0)(747) and tmr_registers(1)(747)) or                                            
                            (tmr_registers(1)(747) and tmr_registers(2)(747)) or                                                       
                            (tmr_registers(0)(747) and tmr_registers(2)(747));                                                         
                                                                                                                                     
        global_tmr_voter(0)(748)  <=    (tmr_registers(0)(748) and tmr_registers(1)(748)) or                                            
                            (tmr_registers(1)(748) and tmr_registers(2)(748)) or                                                       
                            (tmr_registers(0)(748) and tmr_registers(2)(748));                                                         
                                                                                                                                     
        global_tmr_voter(0)(749)  <=    (tmr_registers(0)(749) and tmr_registers(1)(749)) or                                            
                            (tmr_registers(1)(749) and tmr_registers(2)(749)) or                                                       
                            (tmr_registers(0)(749) and tmr_registers(2)(749));                                                         
                                                                                                                                     
        global_tmr_voter(0)(750)  <=    (tmr_registers(0)(750) and tmr_registers(1)(750)) or                                            
                            (tmr_registers(1)(750) and tmr_registers(2)(750)) or                                                       
                            (tmr_registers(0)(750) and tmr_registers(2)(750));                                                         
                                                                                                                                     
        global_tmr_voter(0)(751)  <=    (tmr_registers(0)(751) and tmr_registers(1)(751)) or                                            
                            (tmr_registers(1)(751) and tmr_registers(2)(751)) or                                                       
                            (tmr_registers(0)(751) and tmr_registers(2)(751));                                                         
                                                                                                                                     
        global_tmr_voter(0)(752)  <=    (tmr_registers(0)(752) and tmr_registers(1)(752)) or                                            
                            (tmr_registers(1)(752) and tmr_registers(2)(752)) or                                                       
                            (tmr_registers(0)(752) and tmr_registers(2)(752));                                                         
                                                                                                                                     
        global_tmr_voter(0)(753)  <=    (tmr_registers(0)(753) and tmr_registers(1)(753)) or                                            
                            (tmr_registers(1)(753) and tmr_registers(2)(753)) or                                                       
                            (tmr_registers(0)(753) and tmr_registers(2)(753));                                                         
                                                                                                                                     
        global_tmr_voter(0)(754)  <=    (tmr_registers(0)(754) and tmr_registers(1)(754)) or                                            
                            (tmr_registers(1)(754) and tmr_registers(2)(754)) or                                                       
                            (tmr_registers(0)(754) and tmr_registers(2)(754));                                                         
                                                                                                                                     
        global_tmr_voter(0)(755)  <=    (tmr_registers(0)(755) and tmr_registers(1)(755)) or                                            
                            (tmr_registers(1)(755) and tmr_registers(2)(755)) or                                                       
                            (tmr_registers(0)(755) and tmr_registers(2)(755));                                                         
                                                                                                                                     
        global_tmr_voter(0)(756)  <=    (tmr_registers(0)(756) and tmr_registers(1)(756)) or                                            
                            (tmr_registers(1)(756) and tmr_registers(2)(756)) or                                                       
                            (tmr_registers(0)(756) and tmr_registers(2)(756));                                                         
                                                                                                                                     
        global_tmr_voter(0)(757)  <=    (tmr_registers(0)(757) and tmr_registers(1)(757)) or                                            
                            (tmr_registers(1)(757) and tmr_registers(2)(757)) or                                                       
                            (tmr_registers(0)(757) and tmr_registers(2)(757));                                                         
                                                                                                                                     
        global_tmr_voter(0)(758)  <=    (tmr_registers(0)(758) and tmr_registers(1)(758)) or                                            
                            (tmr_registers(1)(758) and tmr_registers(2)(758)) or                                                       
                            (tmr_registers(0)(758) and tmr_registers(2)(758));                                                         
                                                                                                                                     
        global_tmr_voter(0)(759)  <=    (tmr_registers(0)(759) and tmr_registers(1)(759)) or                                            
                            (tmr_registers(1)(759) and tmr_registers(2)(759)) or                                                       
                            (tmr_registers(0)(759) and tmr_registers(2)(759));                                                         
                                                                                                                                     
        global_tmr_voter(0)(760)  <=    (tmr_registers(0)(760) and tmr_registers(1)(760)) or                                            
                            (tmr_registers(1)(760) and tmr_registers(2)(760)) or                                                       
                            (tmr_registers(0)(760) and tmr_registers(2)(760));                                                         
                                                                                                                                     
        global_tmr_voter(0)(761)  <=    (tmr_registers(0)(761) and tmr_registers(1)(761)) or                                            
                            (tmr_registers(1)(761) and tmr_registers(2)(761)) or                                                       
                            (tmr_registers(0)(761) and tmr_registers(2)(761));                                                         
                                                                                                                                     
        global_tmr_voter(0)(762)  <=    (tmr_registers(0)(762) and tmr_registers(1)(762)) or                                            
                            (tmr_registers(1)(762) and tmr_registers(2)(762)) or                                                       
                            (tmr_registers(0)(762) and tmr_registers(2)(762));                                                         
                                                                                                                                     
        global_tmr_voter(0)(763)  <=    (tmr_registers(0)(763) and tmr_registers(1)(763)) or                                            
                            (tmr_registers(1)(763) and tmr_registers(2)(763)) or                                                       
                            (tmr_registers(0)(763) and tmr_registers(2)(763));                                                         
                                                                                                                                     
        global_tmr_voter(0)(764)  <=    (tmr_registers(0)(764) and tmr_registers(1)(764)) or                                            
                            (tmr_registers(1)(764) and tmr_registers(2)(764)) or                                                       
                            (tmr_registers(0)(764) and tmr_registers(2)(764));                                                         
                                                                                                                                     
        global_tmr_voter(0)(765)  <=    (tmr_registers(0)(765) and tmr_registers(1)(765)) or                                            
                            (tmr_registers(1)(765) and tmr_registers(2)(765)) or                                                       
                            (tmr_registers(0)(765) and tmr_registers(2)(765));                                                         
                                                                                                                                     
        global_tmr_voter(0)(766)  <=    (tmr_registers(0)(766) and tmr_registers(1)(766)) or                                            
                            (tmr_registers(1)(766) and tmr_registers(2)(766)) or                                                       
                            (tmr_registers(0)(766) and tmr_registers(2)(766));                                                         
                                                                                                                                     
        global_tmr_voter(0)(767)  <=    (tmr_registers(0)(767) and tmr_registers(1)(767)) or                                            
                            (tmr_registers(1)(767) and tmr_registers(2)(767)) or                                                       
                            (tmr_registers(0)(767) and tmr_registers(2)(767));                                                         
                                                                                                                                     
        global_tmr_voter(0)(768)  <=    (tmr_registers(0)(768) and tmr_registers(1)(768)) or                                            
                            (tmr_registers(1)(768) and tmr_registers(2)(768)) or                                                       
                            (tmr_registers(0)(768) and tmr_registers(2)(768));                                                         
                                                                                                                                     
        global_tmr_voter(0)(769)  <=    (tmr_registers(0)(769) and tmr_registers(1)(769)) or                                            
                            (tmr_registers(1)(769) and tmr_registers(2)(769)) or                                                       
                            (tmr_registers(0)(769) and tmr_registers(2)(769));                                                         
                                                                                                                                     
        global_tmr_voter(0)(770)  <=    (tmr_registers(0)(770) and tmr_registers(1)(770)) or                                            
                            (tmr_registers(1)(770) and tmr_registers(2)(770)) or                                                       
                            (tmr_registers(0)(770) and tmr_registers(2)(770));                                                         
                                                                                                                                     
        global_tmr_voter(0)(771)  <=    (tmr_registers(0)(771) and tmr_registers(1)(771)) or                                            
                            (tmr_registers(1)(771) and tmr_registers(2)(771)) or                                                       
                            (tmr_registers(0)(771) and tmr_registers(2)(771));                                                         
                                                                                                                                     
        global_tmr_voter(0)(772)  <=    (tmr_registers(0)(772) and tmr_registers(1)(772)) or                                            
                            (tmr_registers(1)(772) and tmr_registers(2)(772)) or                                                       
                            (tmr_registers(0)(772) and tmr_registers(2)(772));                                                         
                                                                                                                                     
        global_tmr_voter(0)(773)  <=    (tmr_registers(0)(773) and tmr_registers(1)(773)) or                                            
                            (tmr_registers(1)(773) and tmr_registers(2)(773)) or                                                       
                            (tmr_registers(0)(773) and tmr_registers(2)(773));                                                         
                                                                                                                                     
        global_tmr_voter(0)(774)  <=    (tmr_registers(0)(774) and tmr_registers(1)(774)) or                                            
                            (tmr_registers(1)(774) and tmr_registers(2)(774)) or                                                       
                            (tmr_registers(0)(774) and tmr_registers(2)(774));                                                         
                                                                                                                                     
        global_tmr_voter(0)(775)  <=    (tmr_registers(0)(775) and tmr_registers(1)(775)) or                                            
                            (tmr_registers(1)(775) and tmr_registers(2)(775)) or                                                       
                            (tmr_registers(0)(775) and tmr_registers(2)(775));                                                         
                                                                                                                                     
        global_tmr_voter(0)(776)  <=    (tmr_registers(0)(776) and tmr_registers(1)(776)) or                                            
                            (tmr_registers(1)(776) and tmr_registers(2)(776)) or                                                       
                            (tmr_registers(0)(776) and tmr_registers(2)(776));                                                         
                                                                                                                                     
        global_tmr_voter(0)(777)  <=    (tmr_registers(0)(777) and tmr_registers(1)(777)) or                                            
                            (tmr_registers(1)(777) and tmr_registers(2)(777)) or                                                       
                            (tmr_registers(0)(777) and tmr_registers(2)(777));                                                         
                                                                                                                                     
        global_tmr_voter(0)(778)  <=    (tmr_registers(0)(778) and tmr_registers(1)(778)) or                                            
                            (tmr_registers(1)(778) and tmr_registers(2)(778)) or                                                       
                            (tmr_registers(0)(778) and tmr_registers(2)(778));                                                         
                                                                                                                                     
        global_tmr_voter(0)(779)  <=    (tmr_registers(0)(779) and tmr_registers(1)(779)) or                                            
                            (tmr_registers(1)(779) and tmr_registers(2)(779)) or                                                       
                            (tmr_registers(0)(779) and tmr_registers(2)(779));                                                         
                                                                                                                                     
        global_tmr_voter(0)(780)  <=    (tmr_registers(0)(780) and tmr_registers(1)(780)) or                                            
                            (tmr_registers(1)(780) and tmr_registers(2)(780)) or                                                       
                            (tmr_registers(0)(780) and tmr_registers(2)(780));                                                         
                                                                                                                                     
        global_tmr_voter(0)(781)  <=    (tmr_registers(0)(781) and tmr_registers(1)(781)) or                                            
                            (tmr_registers(1)(781) and tmr_registers(2)(781)) or                                                       
                            (tmr_registers(0)(781) and tmr_registers(2)(781));                                                         
                                                                                                                                     
        global_tmr_voter(0)(782)  <=    (tmr_registers(0)(782) and tmr_registers(1)(782)) or                                            
                            (tmr_registers(1)(782) and tmr_registers(2)(782)) or                                                       
                            (tmr_registers(0)(782) and tmr_registers(2)(782));                                                         
                                                                                                                                     
        global_tmr_voter(0)(783)  <=    (tmr_registers(0)(783) and tmr_registers(1)(783)) or                                            
                            (tmr_registers(1)(783) and tmr_registers(2)(783)) or                                                       
                            (tmr_registers(0)(783) and tmr_registers(2)(783));                                                         
                                                                                                                                     
        global_tmr_voter(0)(784)  <=    (tmr_registers(0)(784) and tmr_registers(1)(784)) or                                            
                            (tmr_registers(1)(784) and tmr_registers(2)(784)) or                                                       
                            (tmr_registers(0)(784) and tmr_registers(2)(784));                                                         
                                                                                                                                     
        global_tmr_voter(0)(785)  <=    (tmr_registers(0)(785) and tmr_registers(1)(785)) or                                            
                            (tmr_registers(1)(785) and tmr_registers(2)(785)) or                                                       
                            (tmr_registers(0)(785) and tmr_registers(2)(785));                                                         
                                                                                                                                     
        global_tmr_voter(0)(786)  <=    (tmr_registers(0)(786) and tmr_registers(1)(786)) or                                            
                            (tmr_registers(1)(786) and tmr_registers(2)(786)) or                                                       
                            (tmr_registers(0)(786) and tmr_registers(2)(786));                                                         
                                                                                                                                     
        global_tmr_voter(0)(787)  <=    (tmr_registers(0)(787) and tmr_registers(1)(787)) or                                            
                            (tmr_registers(1)(787) and tmr_registers(2)(787)) or                                                       
                            (tmr_registers(0)(787) and tmr_registers(2)(787));                                                         
                                                                                                                                     
        global_tmr_voter(0)(788)  <=    (tmr_registers(0)(788) and tmr_registers(1)(788)) or                                            
                            (tmr_registers(1)(788) and tmr_registers(2)(788)) or                                                       
                            (tmr_registers(0)(788) and tmr_registers(2)(788));                                                         
                                                                                                                                     
        global_tmr_voter(0)(789)  <=    (tmr_registers(0)(789) and tmr_registers(1)(789)) or                                            
                            (tmr_registers(1)(789) and tmr_registers(2)(789)) or                                                       
                            (tmr_registers(0)(789) and tmr_registers(2)(789));                                                         
                                                                                                                                     
        global_tmr_voter(0)(790)  <=    (tmr_registers(0)(790) and tmr_registers(1)(790)) or                                            
                            (tmr_registers(1)(790) and tmr_registers(2)(790)) or                                                       
                            (tmr_registers(0)(790) and tmr_registers(2)(790));                                                         
                                                                                                                                     
        global_tmr_voter(0)(791)  <=    (tmr_registers(0)(791) and tmr_registers(1)(791)) or                                            
                            (tmr_registers(1)(791) and tmr_registers(2)(791)) or                                                       
                            (tmr_registers(0)(791) and tmr_registers(2)(791));                                                         
                                                                                                                                     
        global_tmr_voter(0)(792)  <=    (tmr_registers(0)(792) and tmr_registers(1)(792)) or                                            
                            (tmr_registers(1)(792) and tmr_registers(2)(792)) or                                                       
                            (tmr_registers(0)(792) and tmr_registers(2)(792));                                                         
                                                                                                                                     
        global_tmr_voter(0)(793)  <=    (tmr_registers(0)(793) and tmr_registers(1)(793)) or                                            
                            (tmr_registers(1)(793) and tmr_registers(2)(793)) or                                                       
                            (tmr_registers(0)(793) and tmr_registers(2)(793));                                                         
                                                                                                                                     
        global_tmr_voter(0)(794)  <=    (tmr_registers(0)(794) and tmr_registers(1)(794)) or                                            
                            (tmr_registers(1)(794) and tmr_registers(2)(794)) or                                                       
                            (tmr_registers(0)(794) and tmr_registers(2)(794));                                                         
                                                                                                                                     
        global_tmr_voter(0)(795)  <=    (tmr_registers(0)(795) and tmr_registers(1)(795)) or                                            
                            (tmr_registers(1)(795) and tmr_registers(2)(795)) or                                                       
                            (tmr_registers(0)(795) and tmr_registers(2)(795));                                                         
                                                                                                                                     
        global_tmr_voter(0)(796)  <=    (tmr_registers(0)(796) and tmr_registers(1)(796)) or                                            
                            (tmr_registers(1)(796) and tmr_registers(2)(796)) or                                                       
                            (tmr_registers(0)(796) and tmr_registers(2)(796));                                                         
                                                                                                                                     
        global_tmr_voter(0)(797)  <=    (tmr_registers(0)(797) and tmr_registers(1)(797)) or                                            
                            (tmr_registers(1)(797) and tmr_registers(2)(797)) or                                                       
                            (tmr_registers(0)(797) and tmr_registers(2)(797));                                                         
                                                                                                                                     
        global_tmr_voter(0)(798)  <=    (tmr_registers(0)(798) and tmr_registers(1)(798)) or                                            
                            (tmr_registers(1)(798) and tmr_registers(2)(798)) or                                                       
                            (tmr_registers(0)(798) and tmr_registers(2)(798));                                                         
                                                                                                                                     
        global_tmr_voter(0)(799)  <=    (tmr_registers(0)(799) and tmr_registers(1)(799)) or                                            
                            (tmr_registers(1)(799) and tmr_registers(2)(799)) or                                                       
                            (tmr_registers(0)(799) and tmr_registers(2)(799));                                                         
                                                                                                                                     
        global_tmr_voter(0)(800)  <=    (tmr_registers(0)(800) and tmr_registers(1)(800)) or                                            
                            (tmr_registers(1)(800) and tmr_registers(2)(800)) or                                                       
                            (tmr_registers(0)(800) and tmr_registers(2)(800));                                                         
                                                                                                                                     
        global_tmr_voter(0)(801)  <=    (tmr_registers(0)(801) and tmr_registers(1)(801)) or                                            
                            (tmr_registers(1)(801) and tmr_registers(2)(801)) or                                                       
                            (tmr_registers(0)(801) and tmr_registers(2)(801));                                                         
                                                                                                                                     
        global_tmr_voter(0)(802)  <=    (tmr_registers(0)(802) and tmr_registers(1)(802)) or                                            
                            (tmr_registers(1)(802) and tmr_registers(2)(802)) or                                                       
                            (tmr_registers(0)(802) and tmr_registers(2)(802));                                                         
                                                                                                                                     
        global_tmr_voter(0)(803)  <=    (tmr_registers(0)(803) and tmr_registers(1)(803)) or                                            
                            (tmr_registers(1)(803) and tmr_registers(2)(803)) or                                                       
                            (tmr_registers(0)(803) and tmr_registers(2)(803));                                                         
                                                                                                                                     
        global_tmr_voter(0)(804)  <=    (tmr_registers(0)(804) and tmr_registers(1)(804)) or                                            
                            (tmr_registers(1)(804) and tmr_registers(2)(804)) or                                                       
                            (tmr_registers(0)(804) and tmr_registers(2)(804));                                                         
                                                                                                                                     
        global_tmr_voter(0)(805)  <=    (tmr_registers(0)(805) and tmr_registers(1)(805)) or                                            
                            (tmr_registers(1)(805) and tmr_registers(2)(805)) or                                                       
                            (tmr_registers(0)(805) and tmr_registers(2)(805));                                                         
                                                                                                                                     
        global_tmr_voter(0)(806)  <=    (tmr_registers(0)(806) and tmr_registers(1)(806)) or                                            
                            (tmr_registers(1)(806) and tmr_registers(2)(806)) or                                                       
                            (tmr_registers(0)(806) and tmr_registers(2)(806));                                                         
                                                                                                                                     
        global_tmr_voter(0)(807)  <=    (tmr_registers(0)(807) and tmr_registers(1)(807)) or                                            
                            (tmr_registers(1)(807) and tmr_registers(2)(807)) or                                                       
                            (tmr_registers(0)(807) and tmr_registers(2)(807));                                                         
                                                                                                                                     
        global_tmr_voter(0)(808)  <=    (tmr_registers(0)(808) and tmr_registers(1)(808)) or                                            
                            (tmr_registers(1)(808) and tmr_registers(2)(808)) or                                                       
                            (tmr_registers(0)(808) and tmr_registers(2)(808));                                                         
                                                                                                                                     
        global_tmr_voter(0)(809)  <=    (tmr_registers(0)(809) and tmr_registers(1)(809)) or                                            
                            (tmr_registers(1)(809) and tmr_registers(2)(809)) or                                                       
                            (tmr_registers(0)(809) and tmr_registers(2)(809));                                                         
                                                                                                                                     
        global_tmr_voter(0)(810)  <=    (tmr_registers(0)(810) and tmr_registers(1)(810)) or                                            
                            (tmr_registers(1)(810) and tmr_registers(2)(810)) or                                                       
                            (tmr_registers(0)(810) and tmr_registers(2)(810));                                                         
                                                                                                                                     
        global_tmr_voter(0)(811)  <=    (tmr_registers(0)(811) and tmr_registers(1)(811)) or                                            
                            (tmr_registers(1)(811) and tmr_registers(2)(811)) or                                                       
                            (tmr_registers(0)(811) and tmr_registers(2)(811));                                                         
                                                                                                                                     
        global_tmr_voter(0)(812)  <=    (tmr_registers(0)(812) and tmr_registers(1)(812)) or                                            
                            (tmr_registers(1)(812) and tmr_registers(2)(812)) or                                                       
                            (tmr_registers(0)(812) and tmr_registers(2)(812));                                                         
                                                                                                                                     
        global_tmr_voter(0)(813)  <=    (tmr_registers(0)(813) and tmr_registers(1)(813)) or                                            
                            (tmr_registers(1)(813) and tmr_registers(2)(813)) or                                                       
                            (tmr_registers(0)(813) and tmr_registers(2)(813));                                                         
                                                                                                                                     
        global_tmr_voter(0)(814)  <=    (tmr_registers(0)(814) and tmr_registers(1)(814)) or                                            
                            (tmr_registers(1)(814) and tmr_registers(2)(814)) or                                                       
                            (tmr_registers(0)(814) and tmr_registers(2)(814));                                                         
                                                                                                                                     
        global_tmr_voter(0)(815)  <=    (tmr_registers(0)(815) and tmr_registers(1)(815)) or                                            
                            (tmr_registers(1)(815) and tmr_registers(2)(815)) or                                                       
                            (tmr_registers(0)(815) and tmr_registers(2)(815));                                                         
                                                                                                                                     
        global_tmr_voter(0)(816)  <=    (tmr_registers(0)(816) and tmr_registers(1)(816)) or                                            
                            (tmr_registers(1)(816) and tmr_registers(2)(816)) or                                                       
                            (tmr_registers(0)(816) and tmr_registers(2)(816));                                                         
                                                                                                                                     
        global_tmr_voter(0)(817)  <=    (tmr_registers(0)(817) and tmr_registers(1)(817)) or                                            
                            (tmr_registers(1)(817) and tmr_registers(2)(817)) or                                                       
                            (tmr_registers(0)(817) and tmr_registers(2)(817));                                                         
                                                                                                                                     
        global_tmr_voter(0)(818)  <=    (tmr_registers(0)(818) and tmr_registers(1)(818)) or                                            
                            (tmr_registers(1)(818) and tmr_registers(2)(818)) or                                                       
                            (tmr_registers(0)(818) and tmr_registers(2)(818));                                                         
                                                                                                                                     
        global_tmr_voter(0)(819)  <=    (tmr_registers(0)(819) and tmr_registers(1)(819)) or                                            
                            (tmr_registers(1)(819) and tmr_registers(2)(819)) or                                                       
                            (tmr_registers(0)(819) and tmr_registers(2)(819));                                                         
                                                                                                                                     
        global_tmr_voter(0)(820)  <=    (tmr_registers(0)(820) and tmr_registers(1)(820)) or                                            
                            (tmr_registers(1)(820) and tmr_registers(2)(820)) or                                                       
                            (tmr_registers(0)(820) and tmr_registers(2)(820));                                                         
                                                                                                                                     
        global_tmr_voter(0)(821)  <=    (tmr_registers(0)(821) and tmr_registers(1)(821)) or                                            
                            (tmr_registers(1)(821) and tmr_registers(2)(821)) or                                                       
                            (tmr_registers(0)(821) and tmr_registers(2)(821));                                                         
                                                                                                                                     
        global_tmr_voter(0)(822)  <=    (tmr_registers(0)(822) and tmr_registers(1)(822)) or                                            
                            (tmr_registers(1)(822) and tmr_registers(2)(822)) or                                                       
                            (tmr_registers(0)(822) and tmr_registers(2)(822));                                                         
                                                                                                                                     
        global_tmr_voter(0)(823)  <=    (tmr_registers(0)(823) and tmr_registers(1)(823)) or                                            
                            (tmr_registers(1)(823) and tmr_registers(2)(823)) or                                                       
                            (tmr_registers(0)(823) and tmr_registers(2)(823));                                                         
                                                                                                                                     
        global_tmr_voter(0)(824)  <=    (tmr_registers(0)(824) and tmr_registers(1)(824)) or                                            
                            (tmr_registers(1)(824) and tmr_registers(2)(824)) or                                                       
                            (tmr_registers(0)(824) and tmr_registers(2)(824));                                                         
                                                                                                                                     
        global_tmr_voter(0)(825)  <=    (tmr_registers(0)(825) and tmr_registers(1)(825)) or                                            
                            (tmr_registers(1)(825) and tmr_registers(2)(825)) or                                                       
                            (tmr_registers(0)(825) and tmr_registers(2)(825));                                                         
                                                                                                                                     
        global_tmr_voter(0)(826)  <=    (tmr_registers(0)(826) and tmr_registers(1)(826)) or                                            
                            (tmr_registers(1)(826) and tmr_registers(2)(826)) or                                                       
                            (tmr_registers(0)(826) and tmr_registers(2)(826));                                                         
                                                                                                                                     
        global_tmr_voter(0)(827)  <=    (tmr_registers(0)(827) and tmr_registers(1)(827)) or                                            
                            (tmr_registers(1)(827) and tmr_registers(2)(827)) or                                                       
                            (tmr_registers(0)(827) and tmr_registers(2)(827));                                                         
                                                                                                                                     
        global_tmr_voter(0)(828)  <=    (tmr_registers(0)(828) and tmr_registers(1)(828)) or                                            
                            (tmr_registers(1)(828) and tmr_registers(2)(828)) or                                                       
                            (tmr_registers(0)(828) and tmr_registers(2)(828));                                                         
                                                                                                                                     
        global_tmr_voter(0)(829)  <=    (tmr_registers(0)(829) and tmr_registers(1)(829)) or                                            
                            (tmr_registers(1)(829) and tmr_registers(2)(829)) or                                                       
                            (tmr_registers(0)(829) and tmr_registers(2)(829));                                                         
                                                                                                                                     
        global_tmr_voter(0)(830)  <=    (tmr_registers(0)(830) and tmr_registers(1)(830)) or                                            
                            (tmr_registers(1)(830) and tmr_registers(2)(830)) or                                                       
                            (tmr_registers(0)(830) and tmr_registers(2)(830));                                                         
                                                                                                                                     
        global_tmr_voter(0)(831)  <=    (tmr_registers(0)(831) and tmr_registers(1)(831)) or                                            
                            (tmr_registers(1)(831) and tmr_registers(2)(831)) or                                                       
                            (tmr_registers(0)(831) and tmr_registers(2)(831));                                                         
                                                                                                                                     
        global_tmr_voter(0)(832)  <=    (tmr_registers(0)(832) and tmr_registers(1)(832)) or                                            
                            (tmr_registers(1)(832) and tmr_registers(2)(832)) or                                                       
                            (tmr_registers(0)(832) and tmr_registers(2)(832));                                                         
                                                                                                                                     
        global_tmr_voter(0)(833)  <=    (tmr_registers(0)(833) and tmr_registers(1)(833)) or                                            
                            (tmr_registers(1)(833) and tmr_registers(2)(833)) or                                                       
                            (tmr_registers(0)(833) and tmr_registers(2)(833));                                                         
                                                                                                                                     
        global_tmr_voter(0)(834)  <=    (tmr_registers(0)(834) and tmr_registers(1)(834)) or                                            
                            (tmr_registers(1)(834) and tmr_registers(2)(834)) or                                                       
                            (tmr_registers(0)(834) and tmr_registers(2)(834));                                                         
                                                                                                                                     
        global_tmr_voter(0)(835)  <=    (tmr_registers(0)(835) and tmr_registers(1)(835)) or                                            
                            (tmr_registers(1)(835) and tmr_registers(2)(835)) or                                                       
                            (tmr_registers(0)(835) and tmr_registers(2)(835));                                                         
                                                                                                                                     
        global_tmr_voter(0)(836)  <=    (tmr_registers(0)(836) and tmr_registers(1)(836)) or                                            
                            (tmr_registers(1)(836) and tmr_registers(2)(836)) or                                                       
                            (tmr_registers(0)(836) and tmr_registers(2)(836));                                                         
                                                                                                                                     
        global_tmr_voter(0)(837)  <=    (tmr_registers(0)(837) and tmr_registers(1)(837)) or                                            
                            (tmr_registers(1)(837) and tmr_registers(2)(837)) or                                                       
                            (tmr_registers(0)(837) and tmr_registers(2)(837));                                                         
                                                                                                                                     
        global_tmr_voter(0)(838)  <=    (tmr_registers(0)(838) and tmr_registers(1)(838)) or                                            
                            (tmr_registers(1)(838) and tmr_registers(2)(838)) or                                                       
                            (tmr_registers(0)(838) and tmr_registers(2)(838));                                                         
                                                                                                                                     
        global_tmr_voter(0)(839)  <=    (tmr_registers(0)(839) and tmr_registers(1)(839)) or                                            
                            (tmr_registers(1)(839) and tmr_registers(2)(839)) or                                                       
                            (tmr_registers(0)(839) and tmr_registers(2)(839));                                                         
                                                                                                                                     
        global_tmr_voter(0)(840)  <=    (tmr_registers(0)(840) and tmr_registers(1)(840)) or                                            
                            (tmr_registers(1)(840) and tmr_registers(2)(840)) or                                                       
                            (tmr_registers(0)(840) and tmr_registers(2)(840));                                                         
                                                                                                                                     
        global_tmr_voter(0)(841)  <=    (tmr_registers(0)(841) and tmr_registers(1)(841)) or                                            
                            (tmr_registers(1)(841) and tmr_registers(2)(841)) or                                                       
                            (tmr_registers(0)(841) and tmr_registers(2)(841));                                                         
                                                                                                                                     
        global_tmr_voter(0)(842)  <=    (tmr_registers(0)(842) and tmr_registers(1)(842)) or                                            
                            (tmr_registers(1)(842) and tmr_registers(2)(842)) or                                                       
                            (tmr_registers(0)(842) and tmr_registers(2)(842));                                                         
                                                                                                                                     
        global_tmr_voter(0)(843)  <=    (tmr_registers(0)(843) and tmr_registers(1)(843)) or                                            
                            (tmr_registers(1)(843) and tmr_registers(2)(843)) or                                                       
                            (tmr_registers(0)(843) and tmr_registers(2)(843));                                                         
                                                                                                                                     
        global_tmr_voter(0)(844)  <=    (tmr_registers(0)(844) and tmr_registers(1)(844)) or                                            
                            (tmr_registers(1)(844) and tmr_registers(2)(844)) or                                                       
                            (tmr_registers(0)(844) and tmr_registers(2)(844));                                                         
                                                                                                                                     
        global_tmr_voter(0)(845)  <=    (tmr_registers(0)(845) and tmr_registers(1)(845)) or                                            
                            (tmr_registers(1)(845) and tmr_registers(2)(845)) or                                                       
                            (tmr_registers(0)(845) and tmr_registers(2)(845));                                                         
                                                                                                                                     
        global_tmr_voter(0)(846)  <=    (tmr_registers(0)(846) and tmr_registers(1)(846)) or                                            
                            (tmr_registers(1)(846) and tmr_registers(2)(846)) or                                                       
                            (tmr_registers(0)(846) and tmr_registers(2)(846));                                                         
                                                                                                                                     
        global_tmr_voter(0)(847)  <=    (tmr_registers(0)(847) and tmr_registers(1)(847)) or                                            
                            (tmr_registers(1)(847) and tmr_registers(2)(847)) or                                                       
                            (tmr_registers(0)(847) and tmr_registers(2)(847));                                                         
                                                                                                                                     
        global_tmr_voter(0)(848)  <=    (tmr_registers(0)(848) and tmr_registers(1)(848)) or                                            
                            (tmr_registers(1)(848) and tmr_registers(2)(848)) or                                                       
                            (tmr_registers(0)(848) and tmr_registers(2)(848));                                                         
                                                                                                                                     
        global_tmr_voter(0)(849)  <=    (tmr_registers(0)(849) and tmr_registers(1)(849)) or                                            
                            (tmr_registers(1)(849) and tmr_registers(2)(849)) or                                                       
                            (tmr_registers(0)(849) and tmr_registers(2)(849));                                                         
                                                                                                                                     
        global_tmr_voter(0)(850)  <=    (tmr_registers(0)(850) and tmr_registers(1)(850)) or                                            
                            (tmr_registers(1)(850) and tmr_registers(2)(850)) or                                                       
                            (tmr_registers(0)(850) and tmr_registers(2)(850));                                                         
                                                                                                                                     
        global_tmr_voter(0)(851)  <=    (tmr_registers(0)(851) and tmr_registers(1)(851)) or                                            
                            (tmr_registers(1)(851) and tmr_registers(2)(851)) or                                                       
                            (tmr_registers(0)(851) and tmr_registers(2)(851));                                                         
                                                                                                                                     
        global_tmr_voter(0)(852)  <=    (tmr_registers(0)(852) and tmr_registers(1)(852)) or                                            
                            (tmr_registers(1)(852) and tmr_registers(2)(852)) or                                                       
                            (tmr_registers(0)(852) and tmr_registers(2)(852));                                                         
                                                                                                                                     
        global_tmr_voter(0)(853)  <=    (tmr_registers(0)(853) and tmr_registers(1)(853)) or                                            
                            (tmr_registers(1)(853) and tmr_registers(2)(853)) or                                                       
                            (tmr_registers(0)(853) and tmr_registers(2)(853));                                                         
                                                                                                                                     
        global_tmr_voter(0)(854)  <=    (tmr_registers(0)(854) and tmr_registers(1)(854)) or                                            
                            (tmr_registers(1)(854) and tmr_registers(2)(854)) or                                                       
                            (tmr_registers(0)(854) and tmr_registers(2)(854));                                                         
                                                                                                                                     
        global_tmr_voter(0)(855)  <=    (tmr_registers(0)(855) and tmr_registers(1)(855)) or                                            
                            (tmr_registers(1)(855) and tmr_registers(2)(855)) or                                                       
                            (tmr_registers(0)(855) and tmr_registers(2)(855));                                                         
                                                                                                                                     
        global_tmr_voter(0)(856)  <=    (tmr_registers(0)(856) and tmr_registers(1)(856)) or                                            
                            (tmr_registers(1)(856) and tmr_registers(2)(856)) or                                                       
                            (tmr_registers(0)(856) and tmr_registers(2)(856));                                                         
                                                                                                                                     
        global_tmr_voter(0)(857)  <=    (tmr_registers(0)(857) and tmr_registers(1)(857)) or                                            
                            (tmr_registers(1)(857) and tmr_registers(2)(857)) or                                                       
                            (tmr_registers(0)(857) and tmr_registers(2)(857));                                                         
                                                                                                                                     
        global_tmr_voter(0)(858)  <=    (tmr_registers(0)(858) and tmr_registers(1)(858)) or                                            
                            (tmr_registers(1)(858) and tmr_registers(2)(858)) or                                                       
                            (tmr_registers(0)(858) and tmr_registers(2)(858));                                                         
                                                                                                                                     
        global_tmr_voter(0)(859)  <=    (tmr_registers(0)(859) and tmr_registers(1)(859)) or                                            
                            (tmr_registers(1)(859) and tmr_registers(2)(859)) or                                                       
                            (tmr_registers(0)(859) and tmr_registers(2)(859));                                                         
                                                                                                                                     
        global_tmr_voter(0)(860)  <=    (tmr_registers(0)(860) and tmr_registers(1)(860)) or                                            
                            (tmr_registers(1)(860) and tmr_registers(2)(860)) or                                                       
                            (tmr_registers(0)(860) and tmr_registers(2)(860));                                                         
                                                                                                                                     
        global_tmr_voter(0)(861)  <=    (tmr_registers(0)(861) and tmr_registers(1)(861)) or                                            
                            (tmr_registers(1)(861) and tmr_registers(2)(861)) or                                                       
                            (tmr_registers(0)(861) and tmr_registers(2)(861));                                                         
                                                                                                                                     
        global_tmr_voter(0)(862)  <=    (tmr_registers(0)(862) and tmr_registers(1)(862)) or                                            
                            (tmr_registers(1)(862) and tmr_registers(2)(862)) or                                                       
                            (tmr_registers(0)(862) and tmr_registers(2)(862));                                                         
                                                                                                                                     
        global_tmr_voter(0)(863)  <=    (tmr_registers(0)(863) and tmr_registers(1)(863)) or                                            
                            (tmr_registers(1)(863) and tmr_registers(2)(863)) or                                                       
                            (tmr_registers(0)(863) and tmr_registers(2)(863));                                                         
                                                                                                                                     
        global_tmr_voter(0)(864)  <=    (tmr_registers(0)(864) and tmr_registers(1)(864)) or                                            
                            (tmr_registers(1)(864) and tmr_registers(2)(864)) or                                                       
                            (tmr_registers(0)(864) and tmr_registers(2)(864));                                                         
                                                                                                                                     
        global_tmr_voter(0)(865)  <=    (tmr_registers(0)(865) and tmr_registers(1)(865)) or                                            
                            (tmr_registers(1)(865) and tmr_registers(2)(865)) or                                                       
                            (tmr_registers(0)(865) and tmr_registers(2)(865));                                                         
                                                                                                                                     
        global_tmr_voter(0)(866)  <=    (tmr_registers(0)(866) and tmr_registers(1)(866)) or                                            
                            (tmr_registers(1)(866) and tmr_registers(2)(866)) or                                                       
                            (tmr_registers(0)(866) and tmr_registers(2)(866));                                                         
                                                                                                                                     
        global_tmr_voter(0)(867)  <=    (tmr_registers(0)(867) and tmr_registers(1)(867)) or                                            
                            (tmr_registers(1)(867) and tmr_registers(2)(867)) or                                                       
                            (tmr_registers(0)(867) and tmr_registers(2)(867));                                                         
                                                                                                                                     
        global_tmr_voter(0)(868)  <=    (tmr_registers(0)(868) and tmr_registers(1)(868)) or                                            
                            (tmr_registers(1)(868) and tmr_registers(2)(868)) or                                                       
                            (tmr_registers(0)(868) and tmr_registers(2)(868));                                                         
                                                                                                                                     
        global_tmr_voter(0)(869)  <=    (tmr_registers(0)(869) and tmr_registers(1)(869)) or                                            
                            (tmr_registers(1)(869) and tmr_registers(2)(869)) or                                                       
                            (tmr_registers(0)(869) and tmr_registers(2)(869));                                                         
                                                                                                                                     
        global_tmr_voter(0)(870)  <=    (tmr_registers(0)(870) and tmr_registers(1)(870)) or                                            
                            (tmr_registers(1)(870) and tmr_registers(2)(870)) or                                                       
                            (tmr_registers(0)(870) and tmr_registers(2)(870));                                                         
                                                                                                                                     
        global_tmr_voter(0)(871)  <=    (tmr_registers(0)(871) and tmr_registers(1)(871)) or                                            
                            (tmr_registers(1)(871) and tmr_registers(2)(871)) or                                                       
                            (tmr_registers(0)(871) and tmr_registers(2)(871));                                                         
                                                                                                                                     
        global_tmr_voter(0)(872)  <=    (tmr_registers(0)(872) and tmr_registers(1)(872)) or                                            
                            (tmr_registers(1)(872) and tmr_registers(2)(872)) or                                                       
                            (tmr_registers(0)(872) and tmr_registers(2)(872));                                                         
                                                                                                                                     
        global_tmr_voter(0)(873)  <=    (tmr_registers(0)(873) and tmr_registers(1)(873)) or                                            
                            (tmr_registers(1)(873) and tmr_registers(2)(873)) or                                                       
                            (tmr_registers(0)(873) and tmr_registers(2)(873));                                                         
                                                                                                                                     
        global_tmr_voter(0)(874)  <=    (tmr_registers(0)(874) and tmr_registers(1)(874)) or                                            
                            (tmr_registers(1)(874) and tmr_registers(2)(874)) or                                                       
                            (tmr_registers(0)(874) and tmr_registers(2)(874));                                                         
                                                                                                                                     
        global_tmr_voter(0)(875)  <=    (tmr_registers(0)(875) and tmr_registers(1)(875)) or                                            
                            (tmr_registers(1)(875) and tmr_registers(2)(875)) or                                                       
                            (tmr_registers(0)(875) and tmr_registers(2)(875));                                                         
                                                                                                                                     
        global_tmr_voter(0)(876)  <=    (tmr_registers(0)(876) and tmr_registers(1)(876)) or                                            
                            (tmr_registers(1)(876) and tmr_registers(2)(876)) or                                                       
                            (tmr_registers(0)(876) and tmr_registers(2)(876));                                                         
                                                                                                                                     
        global_tmr_voter(0)(877)  <=    (tmr_registers(0)(877) and tmr_registers(1)(877)) or                                            
                            (tmr_registers(1)(877) and tmr_registers(2)(877)) or                                                       
                            (tmr_registers(0)(877) and tmr_registers(2)(877));                                                         
                                                                                                                                     
        global_tmr_voter(0)(878)  <=    (tmr_registers(0)(878) and tmr_registers(1)(878)) or                                            
                            (tmr_registers(1)(878) and tmr_registers(2)(878)) or                                                       
                            (tmr_registers(0)(878) and tmr_registers(2)(878));                                                         
                                                                                                                                     
        global_tmr_voter(0)(879)  <=    (tmr_registers(0)(879) and tmr_registers(1)(879)) or                                            
                            (tmr_registers(1)(879) and tmr_registers(2)(879)) or                                                       
                            (tmr_registers(0)(879) and tmr_registers(2)(879));                                                         
                                                                                                                                     
        global_tmr_voter(0)(880)  <=    (tmr_registers(0)(880) and tmr_registers(1)(880)) or                                            
                            (tmr_registers(1)(880) and tmr_registers(2)(880)) or                                                       
                            (tmr_registers(0)(880) and tmr_registers(2)(880));                                                         
                                                                                                                                     
        global_tmr_voter(0)(881)  <=    (tmr_registers(0)(881) and tmr_registers(1)(881)) or                                            
                            (tmr_registers(1)(881) and tmr_registers(2)(881)) or                                                       
                            (tmr_registers(0)(881) and tmr_registers(2)(881));                                                         
                                                                                                                                     
        global_tmr_voter(0)(882)  <=    (tmr_registers(0)(882) and tmr_registers(1)(882)) or                                            
                            (tmr_registers(1)(882) and tmr_registers(2)(882)) or                                                       
                            (tmr_registers(0)(882) and tmr_registers(2)(882));                                                         
                                                                                                                                     
        global_tmr_voter(0)(883)  <=    (tmr_registers(0)(883) and tmr_registers(1)(883)) or                                            
                            (tmr_registers(1)(883) and tmr_registers(2)(883)) or                                                       
                            (tmr_registers(0)(883) and tmr_registers(2)(883));                                                         
                                                                                                                                     
        global_tmr_voter(0)(884)  <=    (tmr_registers(0)(884) and tmr_registers(1)(884)) or                                            
                            (tmr_registers(1)(884) and tmr_registers(2)(884)) or                                                       
                            (tmr_registers(0)(884) and tmr_registers(2)(884));                                                         
                                                                                                                                     
        global_tmr_voter(0)(885)  <=    (tmr_registers(0)(885) and tmr_registers(1)(885)) or                                            
                            (tmr_registers(1)(885) and tmr_registers(2)(885)) or                                                       
                            (tmr_registers(0)(885) and tmr_registers(2)(885));                                                         
                                                                                                                                     
        global_tmr_voter(0)(886)  <=    (tmr_registers(0)(886) and tmr_registers(1)(886)) or                                            
                            (tmr_registers(1)(886) and tmr_registers(2)(886)) or                                                       
                            (tmr_registers(0)(886) and tmr_registers(2)(886));                                                         
                                                                                                                                     
        global_tmr_voter(0)(887)  <=    (tmr_registers(0)(887) and tmr_registers(1)(887)) or                                            
                            (tmr_registers(1)(887) and tmr_registers(2)(887)) or                                                       
                            (tmr_registers(0)(887) and tmr_registers(2)(887));                                                         
                                                                                                                                     
        global_tmr_voter(0)(888)  <=    (tmr_registers(0)(888) and tmr_registers(1)(888)) or                                            
                            (tmr_registers(1)(888) and tmr_registers(2)(888)) or                                                       
                            (tmr_registers(0)(888) and tmr_registers(2)(888));                                                         
                                                                                                                                     
        global_tmr_voter(0)(889)  <=    (tmr_registers(0)(889) and tmr_registers(1)(889)) or                                            
                            (tmr_registers(1)(889) and tmr_registers(2)(889)) or                                                       
                            (tmr_registers(0)(889) and tmr_registers(2)(889));                                                         
                                                                                                                                     
        global_tmr_voter(0)(890)  <=    (tmr_registers(0)(890) and tmr_registers(1)(890)) or                                            
                            (tmr_registers(1)(890) and tmr_registers(2)(890)) or                                                       
                            (tmr_registers(0)(890) and tmr_registers(2)(890));                                                         
                                                                                                                                     
        global_tmr_voter(0)(891)  <=    (tmr_registers(0)(891) and tmr_registers(1)(891)) or                                            
                            (tmr_registers(1)(891) and tmr_registers(2)(891)) or                                                       
                            (tmr_registers(0)(891) and tmr_registers(2)(891));                                                         
                                                                                                                                     
        global_tmr_voter(0)(892)  <=    (tmr_registers(0)(892) and tmr_registers(1)(892)) or                                            
                            (tmr_registers(1)(892) and tmr_registers(2)(892)) or                                                       
                            (tmr_registers(0)(892) and tmr_registers(2)(892));                                                         
                                                                                                                                     
        global_tmr_voter(0)(893)  <=    (tmr_registers(0)(893) and tmr_registers(1)(893)) or                                            
                            (tmr_registers(1)(893) and tmr_registers(2)(893)) or                                                       
                            (tmr_registers(0)(893) and tmr_registers(2)(893));                                                         
                                                                                                                                     
        global_tmr_voter(0)(894)  <=    (tmr_registers(0)(894) and tmr_registers(1)(894)) or                                            
                            (tmr_registers(1)(894) and tmr_registers(2)(894)) or                                                       
                            (tmr_registers(0)(894) and tmr_registers(2)(894));                                                         
                                                                                                                                     
        global_tmr_voter(0)(895)  <=    (tmr_registers(0)(895) and tmr_registers(1)(895)) or                                            
                            (tmr_registers(1)(895) and tmr_registers(2)(895)) or                                                       
                            (tmr_registers(0)(895) and tmr_registers(2)(895));                                                         
                                                                                                                                     
        global_tmr_voter(0)(896)  <=    (tmr_registers(0)(896) and tmr_registers(1)(896)) or                                            
                            (tmr_registers(1)(896) and tmr_registers(2)(896)) or                                                       
                            (tmr_registers(0)(896) and tmr_registers(2)(896));                                                         
                                                                                                                                     
        global_tmr_voter(0)(897)  <=    (tmr_registers(0)(897) and tmr_registers(1)(897)) or                                            
                            (tmr_registers(1)(897) and tmr_registers(2)(897)) or                                                       
                            (tmr_registers(0)(897) and tmr_registers(2)(897));                                                         
                                                                                                                                     
        global_tmr_voter(0)(898)  <=    (tmr_registers(0)(898) and tmr_registers(1)(898)) or                                            
                            (tmr_registers(1)(898) and tmr_registers(2)(898)) or                                                       
                            (tmr_registers(0)(898) and tmr_registers(2)(898));                                                         
                                                                                                                                     
        global_tmr_voter(0)(899)  <=    (tmr_registers(0)(899) and tmr_registers(1)(899)) or                                            
                            (tmr_registers(1)(899) and tmr_registers(2)(899)) or                                                       
                            (tmr_registers(0)(899) and tmr_registers(2)(899));                                                         
                                                                                                                                     
        global_tmr_voter(0)(900)  <=    (tmr_registers(0)(900) and tmr_registers(1)(900)) or                                            
                            (tmr_registers(1)(900) and tmr_registers(2)(900)) or                                                       
                            (tmr_registers(0)(900) and tmr_registers(2)(900));                                                         
                                                                                                                                     
        global_tmr_voter(0)(901)  <=    (tmr_registers(0)(901) and tmr_registers(1)(901)) or                                            
                            (tmr_registers(1)(901) and tmr_registers(2)(901)) or                                                       
                            (tmr_registers(0)(901) and tmr_registers(2)(901));                                                         
                                                                                                                                     
        global_tmr_voter(0)(902)  <=    (tmr_registers(0)(902) and tmr_registers(1)(902)) or                                            
                            (tmr_registers(1)(902) and tmr_registers(2)(902)) or                                                       
                            (tmr_registers(0)(902) and tmr_registers(2)(902));                                                         
                                                                                                                                     
        global_tmr_voter(0)(903)  <=    (tmr_registers(0)(903) and tmr_registers(1)(903)) or                                            
                            (tmr_registers(1)(903) and tmr_registers(2)(903)) or                                                       
                            (tmr_registers(0)(903) and tmr_registers(2)(903));                                                         
                                                                                                                                     
        global_tmr_voter(0)(904)  <=    (tmr_registers(0)(904) and tmr_registers(1)(904)) or                                            
                            (tmr_registers(1)(904) and tmr_registers(2)(904)) or                                                       
                            (tmr_registers(0)(904) and tmr_registers(2)(904));                                                         
                                                                                                                                     
        global_tmr_voter(0)(905)  <=    (tmr_registers(0)(905) and tmr_registers(1)(905)) or                                            
                            (tmr_registers(1)(905) and tmr_registers(2)(905)) or                                                       
                            (tmr_registers(0)(905) and tmr_registers(2)(905));                                                         
                                                                                                                                     
        global_tmr_voter(0)(906)  <=    (tmr_registers(0)(906) and tmr_registers(1)(906)) or                                            
                            (tmr_registers(1)(906) and tmr_registers(2)(906)) or                                                       
                            (tmr_registers(0)(906) and tmr_registers(2)(906));                                                         
                                                                                                                                     
        global_tmr_voter(0)(907)  <=    (tmr_registers(0)(907) and tmr_registers(1)(907)) or                                            
                            (tmr_registers(1)(907) and tmr_registers(2)(907)) or                                                       
                            (tmr_registers(0)(907) and tmr_registers(2)(907));                                                         
                                                                                                                                     
        global_tmr_voter(0)(908)  <=    (tmr_registers(0)(908) and tmr_registers(1)(908)) or                                            
                            (tmr_registers(1)(908) and tmr_registers(2)(908)) or                                                       
                            (tmr_registers(0)(908) and tmr_registers(2)(908));                                                         
                                                                                                                                     
        global_tmr_voter(0)(909)  <=    (tmr_registers(0)(909) and tmr_registers(1)(909)) or                                            
                            (tmr_registers(1)(909) and tmr_registers(2)(909)) or                                                       
                            (tmr_registers(0)(909) and tmr_registers(2)(909));                                                         
                                                                                                                                     
        global_tmr_voter(0)(910)  <=    (tmr_registers(0)(910) and tmr_registers(1)(910)) or                                            
                            (tmr_registers(1)(910) and tmr_registers(2)(910)) or                                                       
                            (tmr_registers(0)(910) and tmr_registers(2)(910));                                                         
                                                                                                                                     
        global_tmr_voter(0)(911)  <=    (tmr_registers(0)(911) and tmr_registers(1)(911)) or                                            
                            (tmr_registers(1)(911) and tmr_registers(2)(911)) or                                                       
                            (tmr_registers(0)(911) and tmr_registers(2)(911));                                                         
                                                                                                                                     
        global_tmr_voter(0)(912)  <=    (tmr_registers(0)(912) and tmr_registers(1)(912)) or                                            
                            (tmr_registers(1)(912) and tmr_registers(2)(912)) or                                                       
                            (tmr_registers(0)(912) and tmr_registers(2)(912));                                                         
                                                                                                                                     
        global_tmr_voter(0)(913)  <=    (tmr_registers(0)(913) and tmr_registers(1)(913)) or                                            
                            (tmr_registers(1)(913) and tmr_registers(2)(913)) or                                                       
                            (tmr_registers(0)(913) and tmr_registers(2)(913));                                                         
                                                                                                                                     
        global_tmr_voter(0)(914)  <=    (tmr_registers(0)(914) and tmr_registers(1)(914)) or                                            
                            (tmr_registers(1)(914) and tmr_registers(2)(914)) or                                                       
                            (tmr_registers(0)(914) and tmr_registers(2)(914));                                                         
                                                                                                                                     
        global_tmr_voter(0)(915)  <=    (tmr_registers(0)(915) and tmr_registers(1)(915)) or                                            
                            (tmr_registers(1)(915) and tmr_registers(2)(915)) or                                                       
                            (tmr_registers(0)(915) and tmr_registers(2)(915));                                                         
                                                                                                                                     
        global_tmr_voter(0)(916)  <=    (tmr_registers(0)(916) and tmr_registers(1)(916)) or                                            
                            (tmr_registers(1)(916) and tmr_registers(2)(916)) or                                                       
                            (tmr_registers(0)(916) and tmr_registers(2)(916));                                                         
                                                                                                                                     
        global_tmr_voter(0)(917)  <=    (tmr_registers(0)(917) and tmr_registers(1)(917)) or                                            
                            (tmr_registers(1)(917) and tmr_registers(2)(917)) or                                                       
                            (tmr_registers(0)(917) and tmr_registers(2)(917));                                                         
                                                                                                                                     
        global_tmr_voter(0)(918)  <=    (tmr_registers(0)(918) and tmr_registers(1)(918)) or                                            
                            (tmr_registers(1)(918) and tmr_registers(2)(918)) or                                                       
                            (tmr_registers(0)(918) and tmr_registers(2)(918));                                                         
                                                                                                                                     
        global_tmr_voter(0)(919)  <=    (tmr_registers(0)(919) and tmr_registers(1)(919)) or                                            
                            (tmr_registers(1)(919) and tmr_registers(2)(919)) or                                                       
                            (tmr_registers(0)(919) and tmr_registers(2)(919));                                                         
                                                                                                                                     
        global_tmr_voter(0)(920)  <=    (tmr_registers(0)(920) and tmr_registers(1)(920)) or                                            
                            (tmr_registers(1)(920) and tmr_registers(2)(920)) or                                                       
                            (tmr_registers(0)(920) and tmr_registers(2)(920));                                                         
                                                                                                                                     
        global_tmr_voter(0)(921)  <=    (tmr_registers(0)(921) and tmr_registers(1)(921)) or                                            
                            (tmr_registers(1)(921) and tmr_registers(2)(921)) or                                                       
                            (tmr_registers(0)(921) and tmr_registers(2)(921));                                                         
                                                                                                                                     
        global_tmr_voter(0)(922)  <=    (tmr_registers(0)(922) and tmr_registers(1)(922)) or                                            
                            (tmr_registers(1)(922) and tmr_registers(2)(922)) or                                                       
                            (tmr_registers(0)(922) and tmr_registers(2)(922));                                                         
                                                                                                                                     
        global_tmr_voter(0)(923)  <=    (tmr_registers(0)(923) and tmr_registers(1)(923)) or                                            
                            (tmr_registers(1)(923) and tmr_registers(2)(923)) or                                                       
                            (tmr_registers(0)(923) and tmr_registers(2)(923));                                                         
                                                                                                                                     
        global_tmr_voter(0)(924)  <=    (tmr_registers(0)(924) and tmr_registers(1)(924)) or                                            
                            (tmr_registers(1)(924) and tmr_registers(2)(924)) or                                                       
                            (tmr_registers(0)(924) and tmr_registers(2)(924));                                                         
                                                                                                                                     
        global_tmr_voter(0)(925)  <=    (tmr_registers(0)(925) and tmr_registers(1)(925)) or                                            
                            (tmr_registers(1)(925) and tmr_registers(2)(925)) or                                                       
                            (tmr_registers(0)(925) and tmr_registers(2)(925));                                                         
                                                                                                                                     
        global_tmr_voter(0)(926)  <=    (tmr_registers(0)(926) and tmr_registers(1)(926)) or                                            
                            (tmr_registers(1)(926) and tmr_registers(2)(926)) or                                                       
                            (tmr_registers(0)(926) and tmr_registers(2)(926));                                                         
                                                                                                                                     
        global_tmr_voter(0)(927)  <=    (tmr_registers(0)(927) and tmr_registers(1)(927)) or                                            
                            (tmr_registers(1)(927) and tmr_registers(2)(927)) or                                                       
                            (tmr_registers(0)(927) and tmr_registers(2)(927));                                                         
                                                                                                                                     
        global_tmr_voter(0)(928)  <=    (tmr_registers(0)(928) and tmr_registers(1)(928)) or                                            
                            (tmr_registers(1)(928) and tmr_registers(2)(928)) or                                                       
                            (tmr_registers(0)(928) and tmr_registers(2)(928));                                                         
                                                                                                                                     
        global_tmr_voter(0)(929)  <=    (tmr_registers(0)(929) and tmr_registers(1)(929)) or                                            
                            (tmr_registers(1)(929) and tmr_registers(2)(929)) or                                                       
                            (tmr_registers(0)(929) and tmr_registers(2)(929));                                                         
                                                                                                                                     
        global_tmr_voter(0)(930)  <=    (tmr_registers(0)(930) and tmr_registers(1)(930)) or                                            
                            (tmr_registers(1)(930) and tmr_registers(2)(930)) or                                                       
                            (tmr_registers(0)(930) and tmr_registers(2)(930));                                                         
                                                                                                                                     
        global_tmr_voter(0)(931)  <=    (tmr_registers(0)(931) and tmr_registers(1)(931)) or                                            
                            (tmr_registers(1)(931) and tmr_registers(2)(931)) or                                                       
                            (tmr_registers(0)(931) and tmr_registers(2)(931));                                                         
                                                                                                                                     
        global_tmr_voter(0)(932)  <=    (tmr_registers(0)(932) and tmr_registers(1)(932)) or                                            
                            (tmr_registers(1)(932) and tmr_registers(2)(932)) or                                                       
                            (tmr_registers(0)(932) and tmr_registers(2)(932));                                                         
                                                                                                                                     
        global_tmr_voter(0)(933)  <=    (tmr_registers(0)(933) and tmr_registers(1)(933)) or                                            
                            (tmr_registers(1)(933) and tmr_registers(2)(933)) or                                                       
                            (tmr_registers(0)(933) and tmr_registers(2)(933));                                                         
                                                                                                                                     
        global_tmr_voter(0)(934)  <=    (tmr_registers(0)(934) and tmr_registers(1)(934)) or                                            
                            (tmr_registers(1)(934) and tmr_registers(2)(934)) or                                                       
                            (tmr_registers(0)(934) and tmr_registers(2)(934));                                                         
                                                                                                                                     
        global_tmr_voter(0)(935)  <=    (tmr_registers(0)(935) and tmr_registers(1)(935)) or                                            
                            (tmr_registers(1)(935) and tmr_registers(2)(935)) or                                                       
                            (tmr_registers(0)(935) and tmr_registers(2)(935));                                                         
                                                                                                                                     
        global_tmr_voter(0)(936)  <=    (tmr_registers(0)(936) and tmr_registers(1)(936)) or                                            
                            (tmr_registers(1)(936) and tmr_registers(2)(936)) or                                                       
                            (tmr_registers(0)(936) and tmr_registers(2)(936));                                                         
                                                                                                                                     
        global_tmr_voter(0)(937)  <=    (tmr_registers(0)(937) and tmr_registers(1)(937)) or                                            
                            (tmr_registers(1)(937) and tmr_registers(2)(937)) or                                                       
                            (tmr_registers(0)(937) and tmr_registers(2)(937));                                                         
                                                                                                                                     
        global_tmr_voter(0)(938)  <=    (tmr_registers(0)(938) and tmr_registers(1)(938)) or                                            
                            (tmr_registers(1)(938) and tmr_registers(2)(938)) or                                                       
                            (tmr_registers(0)(938) and tmr_registers(2)(938));                                                         
                                                                                                                                     
        global_tmr_voter(0)(939)  <=    (tmr_registers(0)(939) and tmr_registers(1)(939)) or                                            
                            (tmr_registers(1)(939) and tmr_registers(2)(939)) or                                                       
                            (tmr_registers(0)(939) and tmr_registers(2)(939));                                                         
                                                                                                                                     
        global_tmr_voter(0)(940)  <=    (tmr_registers(0)(940) and tmr_registers(1)(940)) or                                            
                            (tmr_registers(1)(940) and tmr_registers(2)(940)) or                                                       
                            (tmr_registers(0)(940) and tmr_registers(2)(940));                                                         
                                                                                                                                     
        global_tmr_voter(0)(941)  <=    (tmr_registers(0)(941) and tmr_registers(1)(941)) or                                            
                            (tmr_registers(1)(941) and tmr_registers(2)(941)) or                                                       
                            (tmr_registers(0)(941) and tmr_registers(2)(941));                                                         
                                                                                                                                     
        global_tmr_voter(0)(942)  <=    (tmr_registers(0)(942) and tmr_registers(1)(942)) or                                            
                            (tmr_registers(1)(942) and tmr_registers(2)(942)) or                                                       
                            (tmr_registers(0)(942) and tmr_registers(2)(942));                                                         
                                                                                                                                     
        global_tmr_voter(0)(943)  <=    (tmr_registers(0)(943) and tmr_registers(1)(943)) or                                            
                            (tmr_registers(1)(943) and tmr_registers(2)(943)) or                                                       
                            (tmr_registers(0)(943) and tmr_registers(2)(943));                                                         
                                                                                                                                     
        global_tmr_voter(0)(944)  <=    (tmr_registers(0)(944) and tmr_registers(1)(944)) or                                            
                            (tmr_registers(1)(944) and tmr_registers(2)(944)) or                                                       
                            (tmr_registers(0)(944) and tmr_registers(2)(944));                                                         
                                                                                                                                     
        global_tmr_voter(0)(945)  <=    (tmr_registers(0)(945) and tmr_registers(1)(945)) or                                            
                            (tmr_registers(1)(945) and tmr_registers(2)(945)) or                                                       
                            (tmr_registers(0)(945) and tmr_registers(2)(945));                                                         
                                                                                                                                     
        global_tmr_voter(0)(946)  <=    (tmr_registers(0)(946) and tmr_registers(1)(946)) or                                            
                            (tmr_registers(1)(946) and tmr_registers(2)(946)) or                                                       
                            (tmr_registers(0)(946) and tmr_registers(2)(946));                                                         
                                                                                                                                     
        global_tmr_voter(0)(947)  <=    (tmr_registers(0)(947) and tmr_registers(1)(947)) or                                            
                            (tmr_registers(1)(947) and tmr_registers(2)(947)) or                                                       
                            (tmr_registers(0)(947) and tmr_registers(2)(947));                                                         
                                                                                                                                     
        global_tmr_voter(0)(948)  <=    (tmr_registers(0)(948) and tmr_registers(1)(948)) or                                            
                            (tmr_registers(1)(948) and tmr_registers(2)(948)) or                                                       
                            (tmr_registers(0)(948) and tmr_registers(2)(948));                                                         
                                                                                                                                     
        global_tmr_voter(0)(949)  <=    (tmr_registers(0)(949) and tmr_registers(1)(949)) or                                            
                            (tmr_registers(1)(949) and tmr_registers(2)(949)) or                                                       
                            (tmr_registers(0)(949) and tmr_registers(2)(949));                                                         
                                                                                                                                     
        global_tmr_voter(0)(950)  <=    (tmr_registers(0)(950) and tmr_registers(1)(950)) or                                            
                            (tmr_registers(1)(950) and tmr_registers(2)(950)) or                                                       
                            (tmr_registers(0)(950) and tmr_registers(2)(950));                                                         
                                                                                                                                     
        global_tmr_voter(0)(951)  <=    (tmr_registers(0)(951) and tmr_registers(1)(951)) or                                            
                            (tmr_registers(1)(951) and tmr_registers(2)(951)) or                                                       
                            (tmr_registers(0)(951) and tmr_registers(2)(951));                                                         
                                                                                                                                     
        global_tmr_voter(0)(952)  <=    (tmr_registers(0)(952) and tmr_registers(1)(952)) or                                            
                            (tmr_registers(1)(952) and tmr_registers(2)(952)) or                                                       
                            (tmr_registers(0)(952) and tmr_registers(2)(952));                                                         
                                                                                                                                     
        global_tmr_voter(0)(953)  <=    (tmr_registers(0)(953) and tmr_registers(1)(953)) or                                            
                            (tmr_registers(1)(953) and tmr_registers(2)(953)) or                                                       
                            (tmr_registers(0)(953) and tmr_registers(2)(953));                                                         
                                                                                                                                     
        global_tmr_voter(0)(954)  <=    (tmr_registers(0)(954) and tmr_registers(1)(954)) or                                            
                            (tmr_registers(1)(954) and tmr_registers(2)(954)) or                                                       
                            (tmr_registers(0)(954) and tmr_registers(2)(954));                                                         
                                                                                                                                     
        global_tmr_voter(0)(955)  <=    (tmr_registers(0)(955) and tmr_registers(1)(955)) or                                            
                            (tmr_registers(1)(955) and tmr_registers(2)(955)) or                                                       
                            (tmr_registers(0)(955) and tmr_registers(2)(955));                                                         
                                                                                                                                     
        global_tmr_voter(0)(956)  <=    (tmr_registers(0)(956) and tmr_registers(1)(956)) or                                            
                            (tmr_registers(1)(956) and tmr_registers(2)(956)) or                                                       
                            (tmr_registers(0)(956) and tmr_registers(2)(956));                                                         
                                                                                                                                     
        global_tmr_voter(0)(957)  <=    (tmr_registers(0)(957) and tmr_registers(1)(957)) or                                            
                            (tmr_registers(1)(957) and tmr_registers(2)(957)) or                                                       
                            (tmr_registers(0)(957) and tmr_registers(2)(957));                                                         
                                                                                                                                     
        global_tmr_voter(0)(958)  <=    (tmr_registers(0)(958) and tmr_registers(1)(958)) or                                            
                            (tmr_registers(1)(958) and tmr_registers(2)(958)) or                                                       
                            (tmr_registers(0)(958) and tmr_registers(2)(958));                                                         
                                                                                                                                     
        global_tmr_voter(0)(959)  <=    (tmr_registers(0)(959) and tmr_registers(1)(959)) or                                            
                            (tmr_registers(1)(959) and tmr_registers(2)(959)) or                                                       
                            (tmr_registers(0)(959) and tmr_registers(2)(959));                                                         
                                                                                                                                     
        global_tmr_voter(0)(960)  <=    (tmr_registers(0)(960) and tmr_registers(1)(960)) or                                            
                            (tmr_registers(1)(960) and tmr_registers(2)(960)) or                                                       
                            (tmr_registers(0)(960) and tmr_registers(2)(960));                                                         
                                                                                                                                     
        global_tmr_voter(0)(961)  <=    (tmr_registers(0)(961) and tmr_registers(1)(961)) or                                            
                            (tmr_registers(1)(961) and tmr_registers(2)(961)) or                                                       
                            (tmr_registers(0)(961) and tmr_registers(2)(961));                                                         
                                                                                                                                     
        global_tmr_voter(0)(962)  <=    (tmr_registers(0)(962) and tmr_registers(1)(962)) or                                            
                            (tmr_registers(1)(962) and tmr_registers(2)(962)) or                                                       
                            (tmr_registers(0)(962) and tmr_registers(2)(962));                                                         
                                                                                                                                     
        global_tmr_voter(0)(963)  <=    (tmr_registers(0)(963) and tmr_registers(1)(963)) or                                            
                            (tmr_registers(1)(963) and tmr_registers(2)(963)) or                                                       
                            (tmr_registers(0)(963) and tmr_registers(2)(963));                                                         
                                                                                                                                     
        global_tmr_voter(0)(964)  <=    (tmr_registers(0)(964) and tmr_registers(1)(964)) or                                            
                            (tmr_registers(1)(964) and tmr_registers(2)(964)) or                                                       
                            (tmr_registers(0)(964) and tmr_registers(2)(964));                                                         
                                                                                                                                     
        global_tmr_voter(0)(965)  <=    (tmr_registers(0)(965) and tmr_registers(1)(965)) or                                            
                            (tmr_registers(1)(965) and tmr_registers(2)(965)) or                                                       
                            (tmr_registers(0)(965) and tmr_registers(2)(965));                                                         
                                                                                                                                     
        global_tmr_voter(0)(966)  <=    (tmr_registers(0)(966) and tmr_registers(1)(966)) or                                            
                            (tmr_registers(1)(966) and tmr_registers(2)(966)) or                                                       
                            (tmr_registers(0)(966) and tmr_registers(2)(966));                                                         
                                                                                                                                     
        global_tmr_voter(0)(967)  <=    (tmr_registers(0)(967) and tmr_registers(1)(967)) or                                            
                            (tmr_registers(1)(967) and tmr_registers(2)(967)) or                                                       
                            (tmr_registers(0)(967) and tmr_registers(2)(967));                                                         
                                                                                                                                     
        global_tmr_voter(0)(968)  <=    (tmr_registers(0)(968) and tmr_registers(1)(968)) or                                            
                            (tmr_registers(1)(968) and tmr_registers(2)(968)) or                                                       
                            (tmr_registers(0)(968) and tmr_registers(2)(968));                                                         
                                                                                                                                     
        global_tmr_voter(0)(969)  <=    (tmr_registers(0)(969) and tmr_registers(1)(969)) or                                            
                            (tmr_registers(1)(969) and tmr_registers(2)(969)) or                                                       
                            (tmr_registers(0)(969) and tmr_registers(2)(969));                                                         
                                                                                                                                     
        global_tmr_voter(0)(970)  <=    (tmr_registers(0)(970) and tmr_registers(1)(970)) or                                            
                            (tmr_registers(1)(970) and tmr_registers(2)(970)) or                                                       
                            (tmr_registers(0)(970) and tmr_registers(2)(970));                                                         
                                                                                                                                     
        global_tmr_voter(0)(971)  <=    (tmr_registers(0)(971) and tmr_registers(1)(971)) or                                            
                            (tmr_registers(1)(971) and tmr_registers(2)(971)) or                                                       
                            (tmr_registers(0)(971) and tmr_registers(2)(971));                                                         
                                                                                                                                     
        global_tmr_voter(0)(972)  <=    (tmr_registers(0)(972) and tmr_registers(1)(972)) or                                            
                            (tmr_registers(1)(972) and tmr_registers(2)(972)) or                                                       
                            (tmr_registers(0)(972) and tmr_registers(2)(972));                                                         
                                                                                                                                     
        global_tmr_voter(0)(973)  <=    (tmr_registers(0)(973) and tmr_registers(1)(973)) or                                            
                            (tmr_registers(1)(973) and tmr_registers(2)(973)) or                                                       
                            (tmr_registers(0)(973) and tmr_registers(2)(973));                                                         
                                                                                                                                     
        global_tmr_voter(0)(974)  <=    (tmr_registers(0)(974) and tmr_registers(1)(974)) or                                            
                            (tmr_registers(1)(974) and tmr_registers(2)(974)) or                                                       
                            (tmr_registers(0)(974) and tmr_registers(2)(974));                                                         
                                                                                                                                     
        global_tmr_voter(0)(975)  <=    (tmr_registers(0)(975) and tmr_registers(1)(975)) or                                            
                            (tmr_registers(1)(975) and tmr_registers(2)(975)) or                                                       
                            (tmr_registers(0)(975) and tmr_registers(2)(975));                                                         
                                                                                                                                     
        global_tmr_voter(0)(976)  <=    (tmr_registers(0)(976) and tmr_registers(1)(976)) or                                            
                            (tmr_registers(1)(976) and tmr_registers(2)(976)) or                                                       
                            (tmr_registers(0)(976) and tmr_registers(2)(976));                                                         
                                                                                                                                     
        global_tmr_voter(0)(977)  <=    (tmr_registers(0)(977) and tmr_registers(1)(977)) or                                            
                            (tmr_registers(1)(977) and tmr_registers(2)(977)) or                                                       
                            (tmr_registers(0)(977) and tmr_registers(2)(977));                                                         
                                                                                                                                     
        global_tmr_voter(0)(978)  <=    (tmr_registers(0)(978) and tmr_registers(1)(978)) or                                            
                            (tmr_registers(1)(978) and tmr_registers(2)(978)) or                                                       
                            (tmr_registers(0)(978) and tmr_registers(2)(978));                                                         
                                                                                                                                     
        global_tmr_voter(0)(979)  <=    (tmr_registers(0)(979) and tmr_registers(1)(979)) or                                            
                            (tmr_registers(1)(979) and tmr_registers(2)(979)) or                                                       
                            (tmr_registers(0)(979) and tmr_registers(2)(979));                                                         
                                                                                                                                     
        global_tmr_voter(0)(980)  <=    (tmr_registers(0)(980) and tmr_registers(1)(980)) or                                            
                            (tmr_registers(1)(980) and tmr_registers(2)(980)) or                                                       
                            (tmr_registers(0)(980) and tmr_registers(2)(980));                                                         
                                                                                                                                     
        global_tmr_voter(0)(981)  <=    (tmr_registers(0)(981) and tmr_registers(1)(981)) or                                            
                            (tmr_registers(1)(981) and tmr_registers(2)(981)) or                                                       
                            (tmr_registers(0)(981) and tmr_registers(2)(981));                                                         
                                                                                                                                     
        global_tmr_voter(0)(982)  <=    (tmr_registers(0)(982) and tmr_registers(1)(982)) or                                            
                            (tmr_registers(1)(982) and tmr_registers(2)(982)) or                                                       
                            (tmr_registers(0)(982) and tmr_registers(2)(982));                                                         
                                                                                                                                     
        global_tmr_voter(0)(983)  <=    (tmr_registers(0)(983) and tmr_registers(1)(983)) or                                            
                            (tmr_registers(1)(983) and tmr_registers(2)(983)) or                                                       
                            (tmr_registers(0)(983) and tmr_registers(2)(983));                                                         
                                                                                                                                     
        global_tmr_voter(0)(984)  <=    (tmr_registers(0)(984) and tmr_registers(1)(984)) or                                            
                            (tmr_registers(1)(984) and tmr_registers(2)(984)) or                                                       
                            (tmr_registers(0)(984) and tmr_registers(2)(984));                                                         
                                                                                                                                     
        global_tmr_voter(0)(985)  <=    (tmr_registers(0)(985) and tmr_registers(1)(985)) or                                            
                            (tmr_registers(1)(985) and tmr_registers(2)(985)) or                                                       
                            (tmr_registers(0)(985) and tmr_registers(2)(985));                                                         
                                                                                                                                     
        global_tmr_voter(0)(986)  <=    (tmr_registers(0)(986) and tmr_registers(1)(986)) or                                            
                            (tmr_registers(1)(986) and tmr_registers(2)(986)) or                                                       
                            (tmr_registers(0)(986) and tmr_registers(2)(986));                                                         
                                                                                                                                     
        global_tmr_voter(0)(987)  <=    (tmr_registers(0)(987) and tmr_registers(1)(987)) or                                            
                            (tmr_registers(1)(987) and tmr_registers(2)(987)) or                                                       
                            (tmr_registers(0)(987) and tmr_registers(2)(987));                                                         
                                                                                                                                     
        global_tmr_voter(0)(988)  <=    (tmr_registers(0)(988) and tmr_registers(1)(988)) or                                            
                            (tmr_registers(1)(988) and tmr_registers(2)(988)) or                                                       
                            (tmr_registers(0)(988) and tmr_registers(2)(988));                                                         
                                                                                                                                     
        global_tmr_voter(0)(989)  <=    (tmr_registers(0)(989) and tmr_registers(1)(989)) or                                            
                            (tmr_registers(1)(989) and tmr_registers(2)(989)) or                                                       
                            (tmr_registers(0)(989) and tmr_registers(2)(989));                                                         
                                                                                                                                     
        global_tmr_voter(0)(990)  <=    (tmr_registers(0)(990) and tmr_registers(1)(990)) or                                            
                            (tmr_registers(1)(990) and tmr_registers(2)(990)) or                                                       
                            (tmr_registers(0)(990) and tmr_registers(2)(990));                                                         
                                                                                                                                     
        global_tmr_voter(0)(991)  <=    (tmr_registers(0)(991) and tmr_registers(1)(991)) or                                            
                            (tmr_registers(1)(991) and tmr_registers(2)(991)) or                                                       
                            (tmr_registers(0)(991) and tmr_registers(2)(991));                                                         
                                                                                                                                     
        global_tmr_voter(0)(992)  <=    (tmr_registers(0)(992) and tmr_registers(1)(992)) or                                            
                            (tmr_registers(1)(992) and tmr_registers(2)(992)) or                                                       
                            (tmr_registers(0)(992) and tmr_registers(2)(992));                                                         
                                                                                                                                     
        global_tmr_voter(0)(993)  <=    (tmr_registers(0)(993) and tmr_registers(1)(993)) or                                            
                            (tmr_registers(1)(993) and tmr_registers(2)(993)) or                                                       
                            (tmr_registers(0)(993) and tmr_registers(2)(993));                                                         
                                                                                                                                     
        global_tmr_voter(0)(994)  <=    (tmr_registers(0)(994) and tmr_registers(1)(994)) or                                            
                            (tmr_registers(1)(994) and tmr_registers(2)(994)) or                                                       
                            (tmr_registers(0)(994) and tmr_registers(2)(994));                                                         
                                                                                                                                     
        global_tmr_voter(0)(995)  <=    (tmr_registers(0)(995) and tmr_registers(1)(995)) or                                            
                            (tmr_registers(1)(995) and tmr_registers(2)(995)) or                                                       
                            (tmr_registers(0)(995) and tmr_registers(2)(995));                                                         
                                                                                                                                     
        global_tmr_voter(0)(996)  <=    (tmr_registers(0)(996) and tmr_registers(1)(996)) or                                            
                            (tmr_registers(1)(996) and tmr_registers(2)(996)) or                                                       
                            (tmr_registers(0)(996) and tmr_registers(2)(996));                                                         
                                                                                                                                     
        global_tmr_voter(0)(997)  <=    (tmr_registers(0)(997) and tmr_registers(1)(997)) or                                            
                            (tmr_registers(1)(997) and tmr_registers(2)(997)) or                                                       
                            (tmr_registers(0)(997) and tmr_registers(2)(997));                                                         
                                                                                                                                     
        global_tmr_voter(0)(998)  <=    (tmr_registers(0)(998) and tmr_registers(1)(998)) or                                            
                            (tmr_registers(1)(998) and tmr_registers(2)(998)) or                                                       
                            (tmr_registers(0)(998) and tmr_registers(2)(998));                                                         
                                                                                                                                     
        global_tmr_voter(0)(999)  <=    (tmr_registers(0)(999) and tmr_registers(1)(999)) or                                            
                            (tmr_registers(1)(999) and tmr_registers(2)(999)) or                                                       
                            (tmr_registers(0)(999) and tmr_registers(2)(999));                                                         
                                                                                                                                         
                                                                                                                                     
        global_tmr_voter(1)(1)  <=    (tmr_registers(0)(1) and tmr_registers(1)(1)) or                                            
                            (tmr_registers(1)(1) and tmr_registers(2)(1)) or                                                       
                            (tmr_registers(0)(1) and tmr_registers(2)(1));                                                         
                                                                                                                                     
        global_tmr_voter(1)(2)  <=    (tmr_registers(0)(2) and tmr_registers(1)(2)) or                                            
                            (tmr_registers(1)(2) and tmr_registers(2)(2)) or                                                       
                            (tmr_registers(0)(2) and tmr_registers(2)(2));                                                         
                                                                                                                                     
        global_tmr_voter(1)(3)  <=    (tmr_registers(0)(3) and tmr_registers(1)(3)) or                                            
                            (tmr_registers(1)(3) and tmr_registers(2)(3)) or                                                       
                            (tmr_registers(0)(3) and tmr_registers(2)(3));                                                         
                                                                                                                                     
        global_tmr_voter(1)(4)  <=    (tmr_registers(0)(4) and tmr_registers(1)(4)) or                                            
                            (tmr_registers(1)(4) and tmr_registers(2)(4)) or                                                       
                            (tmr_registers(0)(4) and tmr_registers(2)(4));                                                         
                                                                                                                                     
        global_tmr_voter(1)(5)  <=    (tmr_registers(0)(5) and tmr_registers(1)(5)) or                                            
                            (tmr_registers(1)(5) and tmr_registers(2)(5)) or                                                       
                            (tmr_registers(0)(5) and tmr_registers(2)(5));                                                         
                                                                                                                                     
        global_tmr_voter(1)(6)  <=    (tmr_registers(0)(6) and tmr_registers(1)(6)) or                                            
                            (tmr_registers(1)(6) and tmr_registers(2)(6)) or                                                       
                            (tmr_registers(0)(6) and tmr_registers(2)(6));                                                         
                                                                                                                                     
        global_tmr_voter(1)(7)  <=    (tmr_registers(0)(7) and tmr_registers(1)(7)) or                                            
                            (tmr_registers(1)(7) and tmr_registers(2)(7)) or                                                       
                            (tmr_registers(0)(7) and tmr_registers(2)(7));                                                         
                                                                                                                                     
        global_tmr_voter(1)(8)  <=    (tmr_registers(0)(8) and tmr_registers(1)(8)) or                                            
                            (tmr_registers(1)(8) and tmr_registers(2)(8)) or                                                       
                            (tmr_registers(0)(8) and tmr_registers(2)(8));                                                         
                                                                                                                                     
        global_tmr_voter(1)(9)  <=    (tmr_registers(0)(9) and tmr_registers(1)(9)) or                                            
                            (tmr_registers(1)(9) and tmr_registers(2)(9)) or                                                       
                            (tmr_registers(0)(9) and tmr_registers(2)(9));                                                         
                                                                                                                                     
        global_tmr_voter(1)(10)  <=    (tmr_registers(0)(10) and tmr_registers(1)(10)) or                                            
                            (tmr_registers(1)(10) and tmr_registers(2)(10)) or                                                       
                            (tmr_registers(0)(10) and tmr_registers(2)(10));                                                         
                                                                                                                                     
        global_tmr_voter(1)(11)  <=    (tmr_registers(0)(11) and tmr_registers(1)(11)) or                                            
                            (tmr_registers(1)(11) and tmr_registers(2)(11)) or                                                       
                            (tmr_registers(0)(11) and tmr_registers(2)(11));                                                         
                                                                                                                                     
        global_tmr_voter(1)(12)  <=    (tmr_registers(0)(12) and tmr_registers(1)(12)) or                                            
                            (tmr_registers(1)(12) and tmr_registers(2)(12)) or                                                       
                            (tmr_registers(0)(12) and tmr_registers(2)(12));                                                         
                                                                                                                                     
        global_tmr_voter(1)(13)  <=    (tmr_registers(0)(13) and tmr_registers(1)(13)) or                                            
                            (tmr_registers(1)(13) and tmr_registers(2)(13)) or                                                       
                            (tmr_registers(0)(13) and tmr_registers(2)(13));                                                         
                                                                                                                                     
        global_tmr_voter(1)(14)  <=    (tmr_registers(0)(14) and tmr_registers(1)(14)) or                                            
                            (tmr_registers(1)(14) and tmr_registers(2)(14)) or                                                       
                            (tmr_registers(0)(14) and tmr_registers(2)(14));                                                         
                                                                                                                                     
        global_tmr_voter(1)(15)  <=    (tmr_registers(0)(15) and tmr_registers(1)(15)) or                                            
                            (tmr_registers(1)(15) and tmr_registers(2)(15)) or                                                       
                            (tmr_registers(0)(15) and tmr_registers(2)(15));                                                         
                                                                                                                                     
        global_tmr_voter(1)(16)  <=    (tmr_registers(0)(16) and tmr_registers(1)(16)) or                                            
                            (tmr_registers(1)(16) and tmr_registers(2)(16)) or                                                       
                            (tmr_registers(0)(16) and tmr_registers(2)(16));                                                         
                                                                                                                                     
        global_tmr_voter(1)(17)  <=    (tmr_registers(0)(17) and tmr_registers(1)(17)) or                                            
                            (tmr_registers(1)(17) and tmr_registers(2)(17)) or                                                       
                            (tmr_registers(0)(17) and tmr_registers(2)(17));                                                         
                                                                                                                                     
        global_tmr_voter(1)(18)  <=    (tmr_registers(0)(18) and tmr_registers(1)(18)) or                                            
                            (tmr_registers(1)(18) and tmr_registers(2)(18)) or                                                       
                            (tmr_registers(0)(18) and tmr_registers(2)(18));                                                         
                                                                                                                                     
        global_tmr_voter(1)(19)  <=    (tmr_registers(0)(19) and tmr_registers(1)(19)) or                                            
                            (tmr_registers(1)(19) and tmr_registers(2)(19)) or                                                       
                            (tmr_registers(0)(19) and tmr_registers(2)(19));                                                         
                                                                                                                                     
        global_tmr_voter(1)(20)  <=    (tmr_registers(0)(20) and tmr_registers(1)(20)) or                                            
                            (tmr_registers(1)(20) and tmr_registers(2)(20)) or                                                       
                            (tmr_registers(0)(20) and tmr_registers(2)(20));                                                         
                                                                                                                                     
        global_tmr_voter(1)(21)  <=    (tmr_registers(0)(21) and tmr_registers(1)(21)) or                                            
                            (tmr_registers(1)(21) and tmr_registers(2)(21)) or                                                       
                            (tmr_registers(0)(21) and tmr_registers(2)(21));                                                         
                                                                                                                                     
        global_tmr_voter(1)(22)  <=    (tmr_registers(0)(22) and tmr_registers(1)(22)) or                                            
                            (tmr_registers(1)(22) and tmr_registers(2)(22)) or                                                       
                            (tmr_registers(0)(22) and tmr_registers(2)(22));                                                         
                                                                                                                                     
        global_tmr_voter(1)(23)  <=    (tmr_registers(0)(23) and tmr_registers(1)(23)) or                                            
                            (tmr_registers(1)(23) and tmr_registers(2)(23)) or                                                       
                            (tmr_registers(0)(23) and tmr_registers(2)(23));                                                         
                                                                                                                                     
        global_tmr_voter(1)(24)  <=    (tmr_registers(0)(24) and tmr_registers(1)(24)) or                                            
                            (tmr_registers(1)(24) and tmr_registers(2)(24)) or                                                       
                            (tmr_registers(0)(24) and tmr_registers(2)(24));                                                         
                                                                                                                                     
        global_tmr_voter(1)(25)  <=    (tmr_registers(0)(25) and tmr_registers(1)(25)) or                                            
                            (tmr_registers(1)(25) and tmr_registers(2)(25)) or                                                       
                            (tmr_registers(0)(25) and tmr_registers(2)(25));                                                         
                                                                                                                                     
        global_tmr_voter(1)(26)  <=    (tmr_registers(0)(26) and tmr_registers(1)(26)) or                                            
                            (tmr_registers(1)(26) and tmr_registers(2)(26)) or                                                       
                            (tmr_registers(0)(26) and tmr_registers(2)(26));                                                         
                                                                                                                                     
        global_tmr_voter(1)(27)  <=    (tmr_registers(0)(27) and tmr_registers(1)(27)) or                                            
                            (tmr_registers(1)(27) and tmr_registers(2)(27)) or                                                       
                            (tmr_registers(0)(27) and tmr_registers(2)(27));                                                         
                                                                                                                                     
        global_tmr_voter(1)(28)  <=    (tmr_registers(0)(28) and tmr_registers(1)(28)) or                                            
                            (tmr_registers(1)(28) and tmr_registers(2)(28)) or                                                       
                            (tmr_registers(0)(28) and tmr_registers(2)(28));                                                         
                                                                                                                                     
        global_tmr_voter(1)(29)  <=    (tmr_registers(0)(29) and tmr_registers(1)(29)) or                                            
                            (tmr_registers(1)(29) and tmr_registers(2)(29)) or                                                       
                            (tmr_registers(0)(29) and tmr_registers(2)(29));                                                         
                                                                                                                                     
        global_tmr_voter(1)(30)  <=    (tmr_registers(0)(30) and tmr_registers(1)(30)) or                                            
                            (tmr_registers(1)(30) and tmr_registers(2)(30)) or                                                       
                            (tmr_registers(0)(30) and tmr_registers(2)(30));                                                         
                                                                                                                                     
        global_tmr_voter(1)(31)  <=    (tmr_registers(0)(31) and tmr_registers(1)(31)) or                                            
                            (tmr_registers(1)(31) and tmr_registers(2)(31)) or                                                       
                            (tmr_registers(0)(31) and tmr_registers(2)(31));                                                         
                                                                                                                                     
        global_tmr_voter(1)(32)  <=    (tmr_registers(0)(32) and tmr_registers(1)(32)) or                                            
                            (tmr_registers(1)(32) and tmr_registers(2)(32)) or                                                       
                            (tmr_registers(0)(32) and tmr_registers(2)(32));                                                         
                                                                                                                                     
        global_tmr_voter(1)(33)  <=    (tmr_registers(0)(33) and tmr_registers(1)(33)) or                                            
                            (tmr_registers(1)(33) and tmr_registers(2)(33)) or                                                       
                            (tmr_registers(0)(33) and tmr_registers(2)(33));                                                         
                                                                                                                                     
        global_tmr_voter(1)(34)  <=    (tmr_registers(0)(34) and tmr_registers(1)(34)) or                                            
                            (tmr_registers(1)(34) and tmr_registers(2)(34)) or                                                       
                            (tmr_registers(0)(34) and tmr_registers(2)(34));                                                         
                                                                                                                                     
        global_tmr_voter(1)(35)  <=    (tmr_registers(0)(35) and tmr_registers(1)(35)) or                                            
                            (tmr_registers(1)(35) and tmr_registers(2)(35)) or                                                       
                            (tmr_registers(0)(35) and tmr_registers(2)(35));                                                         
                                                                                                                                     
        global_tmr_voter(1)(36)  <=    (tmr_registers(0)(36) and tmr_registers(1)(36)) or                                            
                            (tmr_registers(1)(36) and tmr_registers(2)(36)) or                                                       
                            (tmr_registers(0)(36) and tmr_registers(2)(36));                                                         
                                                                                                                                     
        global_tmr_voter(1)(37)  <=    (tmr_registers(0)(37) and tmr_registers(1)(37)) or                                            
                            (tmr_registers(1)(37) and tmr_registers(2)(37)) or                                                       
                            (tmr_registers(0)(37) and tmr_registers(2)(37));                                                         
                                                                                                                                     
        global_tmr_voter(1)(38)  <=    (tmr_registers(0)(38) and tmr_registers(1)(38)) or                                            
                            (tmr_registers(1)(38) and tmr_registers(2)(38)) or                                                       
                            (tmr_registers(0)(38) and tmr_registers(2)(38));                                                         
                                                                                                                                     
        global_tmr_voter(1)(39)  <=    (tmr_registers(0)(39) and tmr_registers(1)(39)) or                                            
                            (tmr_registers(1)(39) and tmr_registers(2)(39)) or                                                       
                            (tmr_registers(0)(39) and tmr_registers(2)(39));                                                         
                                                                                                                                     
        global_tmr_voter(1)(40)  <=    (tmr_registers(0)(40) and tmr_registers(1)(40)) or                                            
                            (tmr_registers(1)(40) and tmr_registers(2)(40)) or                                                       
                            (tmr_registers(0)(40) and tmr_registers(2)(40));                                                         
                                                                                                                                     
        global_tmr_voter(1)(41)  <=    (tmr_registers(0)(41) and tmr_registers(1)(41)) or                                            
                            (tmr_registers(1)(41) and tmr_registers(2)(41)) or                                                       
                            (tmr_registers(0)(41) and tmr_registers(2)(41));                                                         
                                                                                                                                     
        global_tmr_voter(1)(42)  <=    (tmr_registers(0)(42) and tmr_registers(1)(42)) or                                            
                            (tmr_registers(1)(42) and tmr_registers(2)(42)) or                                                       
                            (tmr_registers(0)(42) and tmr_registers(2)(42));                                                         
                                                                                                                                     
        global_tmr_voter(1)(43)  <=    (tmr_registers(0)(43) and tmr_registers(1)(43)) or                                            
                            (tmr_registers(1)(43) and tmr_registers(2)(43)) or                                                       
                            (tmr_registers(0)(43) and tmr_registers(2)(43));                                                         
                                                                                                                                     
        global_tmr_voter(1)(44)  <=    (tmr_registers(0)(44) and tmr_registers(1)(44)) or                                            
                            (tmr_registers(1)(44) and tmr_registers(2)(44)) or                                                       
                            (tmr_registers(0)(44) and tmr_registers(2)(44));                                                         
                                                                                                                                     
        global_tmr_voter(1)(45)  <=    (tmr_registers(0)(45) and tmr_registers(1)(45)) or                                            
                            (tmr_registers(1)(45) and tmr_registers(2)(45)) or                                                       
                            (tmr_registers(0)(45) and tmr_registers(2)(45));                                                         
                                                                                                                                     
        global_tmr_voter(1)(46)  <=    (tmr_registers(0)(46) and tmr_registers(1)(46)) or                                            
                            (tmr_registers(1)(46) and tmr_registers(2)(46)) or                                                       
                            (tmr_registers(0)(46) and tmr_registers(2)(46));                                                         
                                                                                                                                     
        global_tmr_voter(1)(47)  <=    (tmr_registers(0)(47) and tmr_registers(1)(47)) or                                            
                            (tmr_registers(1)(47) and tmr_registers(2)(47)) or                                                       
                            (tmr_registers(0)(47) and tmr_registers(2)(47));                                                         
                                                                                                                                     
        global_tmr_voter(1)(48)  <=    (tmr_registers(0)(48) and tmr_registers(1)(48)) or                                            
                            (tmr_registers(1)(48) and tmr_registers(2)(48)) or                                                       
                            (tmr_registers(0)(48) and tmr_registers(2)(48));                                                         
                                                                                                                                     
        global_tmr_voter(1)(49)  <=    (tmr_registers(0)(49) and tmr_registers(1)(49)) or                                            
                            (tmr_registers(1)(49) and tmr_registers(2)(49)) or                                                       
                            (tmr_registers(0)(49) and tmr_registers(2)(49));                                                         
                                                                                                                                     
        global_tmr_voter(1)(50)  <=    (tmr_registers(0)(50) and tmr_registers(1)(50)) or                                            
                            (tmr_registers(1)(50) and tmr_registers(2)(50)) or                                                       
                            (tmr_registers(0)(50) and tmr_registers(2)(50));                                                         
                                                                                                                                     
        global_tmr_voter(1)(51)  <=    (tmr_registers(0)(51) and tmr_registers(1)(51)) or                                            
                            (tmr_registers(1)(51) and tmr_registers(2)(51)) or                                                       
                            (tmr_registers(0)(51) and tmr_registers(2)(51));                                                         
                                                                                                                                     
        global_tmr_voter(1)(52)  <=    (tmr_registers(0)(52) and tmr_registers(1)(52)) or                                            
                            (tmr_registers(1)(52) and tmr_registers(2)(52)) or                                                       
                            (tmr_registers(0)(52) and tmr_registers(2)(52));                                                         
                                                                                                                                     
        global_tmr_voter(1)(53)  <=    (tmr_registers(0)(53) and tmr_registers(1)(53)) or                                            
                            (tmr_registers(1)(53) and tmr_registers(2)(53)) or                                                       
                            (tmr_registers(0)(53) and tmr_registers(2)(53));                                                         
                                                                                                                                     
        global_tmr_voter(1)(54)  <=    (tmr_registers(0)(54) and tmr_registers(1)(54)) or                                            
                            (tmr_registers(1)(54) and tmr_registers(2)(54)) or                                                       
                            (tmr_registers(0)(54) and tmr_registers(2)(54));                                                         
                                                                                                                                     
        global_tmr_voter(1)(55)  <=    (tmr_registers(0)(55) and tmr_registers(1)(55)) or                                            
                            (tmr_registers(1)(55) and tmr_registers(2)(55)) or                                                       
                            (tmr_registers(0)(55) and tmr_registers(2)(55));                                                         
                                                                                                                                     
        global_tmr_voter(1)(56)  <=    (tmr_registers(0)(56) and tmr_registers(1)(56)) or                                            
                            (tmr_registers(1)(56) and tmr_registers(2)(56)) or                                                       
                            (tmr_registers(0)(56) and tmr_registers(2)(56));                                                         
                                                                                                                                     
        global_tmr_voter(1)(57)  <=    (tmr_registers(0)(57) and tmr_registers(1)(57)) or                                            
                            (tmr_registers(1)(57) and tmr_registers(2)(57)) or                                                       
                            (tmr_registers(0)(57) and tmr_registers(2)(57));                                                         
                                                                                                                                     
        global_tmr_voter(1)(58)  <=    (tmr_registers(0)(58) and tmr_registers(1)(58)) or                                            
                            (tmr_registers(1)(58) and tmr_registers(2)(58)) or                                                       
                            (tmr_registers(0)(58) and tmr_registers(2)(58));                                                         
                                                                                                                                     
        global_tmr_voter(1)(59)  <=    (tmr_registers(0)(59) and tmr_registers(1)(59)) or                                            
                            (tmr_registers(1)(59) and tmr_registers(2)(59)) or                                                       
                            (tmr_registers(0)(59) and tmr_registers(2)(59));                                                         
                                                                                                                                     
        global_tmr_voter(1)(60)  <=    (tmr_registers(0)(60) and tmr_registers(1)(60)) or                                            
                            (tmr_registers(1)(60) and tmr_registers(2)(60)) or                                                       
                            (tmr_registers(0)(60) and tmr_registers(2)(60));                                                         
                                                                                                                                     
        global_tmr_voter(1)(61)  <=    (tmr_registers(0)(61) and tmr_registers(1)(61)) or                                            
                            (tmr_registers(1)(61) and tmr_registers(2)(61)) or                                                       
                            (tmr_registers(0)(61) and tmr_registers(2)(61));                                                         
                                                                                                                                     
        global_tmr_voter(1)(62)  <=    (tmr_registers(0)(62) and tmr_registers(1)(62)) or                                            
                            (tmr_registers(1)(62) and tmr_registers(2)(62)) or                                                       
                            (tmr_registers(0)(62) and tmr_registers(2)(62));                                                         
                                                                                                                                     
        global_tmr_voter(1)(63)  <=    (tmr_registers(0)(63) and tmr_registers(1)(63)) or                                            
                            (tmr_registers(1)(63) and tmr_registers(2)(63)) or                                                       
                            (tmr_registers(0)(63) and tmr_registers(2)(63));                                                         
                                                                                                                                     
        global_tmr_voter(1)(64)  <=    (tmr_registers(0)(64) and tmr_registers(1)(64)) or                                            
                            (tmr_registers(1)(64) and tmr_registers(2)(64)) or                                                       
                            (tmr_registers(0)(64) and tmr_registers(2)(64));                                                         
                                                                                                                                     
        global_tmr_voter(1)(65)  <=    (tmr_registers(0)(65) and tmr_registers(1)(65)) or                                            
                            (tmr_registers(1)(65) and tmr_registers(2)(65)) or                                                       
                            (tmr_registers(0)(65) and tmr_registers(2)(65));                                                         
                                                                                                                                     
        global_tmr_voter(1)(66)  <=    (tmr_registers(0)(66) and tmr_registers(1)(66)) or                                            
                            (tmr_registers(1)(66) and tmr_registers(2)(66)) or                                                       
                            (tmr_registers(0)(66) and tmr_registers(2)(66));                                                         
                                                                                                                                     
        global_tmr_voter(1)(67)  <=    (tmr_registers(0)(67) and tmr_registers(1)(67)) or                                            
                            (tmr_registers(1)(67) and tmr_registers(2)(67)) or                                                       
                            (tmr_registers(0)(67) and tmr_registers(2)(67));                                                         
                                                                                                                                     
        global_tmr_voter(1)(68)  <=    (tmr_registers(0)(68) and tmr_registers(1)(68)) or                                            
                            (tmr_registers(1)(68) and tmr_registers(2)(68)) or                                                       
                            (tmr_registers(0)(68) and tmr_registers(2)(68));                                                         
                                                                                                                                     
        global_tmr_voter(1)(69)  <=    (tmr_registers(0)(69) and tmr_registers(1)(69)) or                                            
                            (tmr_registers(1)(69) and tmr_registers(2)(69)) or                                                       
                            (tmr_registers(0)(69) and tmr_registers(2)(69));                                                         
                                                                                                                                     
        global_tmr_voter(1)(70)  <=    (tmr_registers(0)(70) and tmr_registers(1)(70)) or                                            
                            (tmr_registers(1)(70) and tmr_registers(2)(70)) or                                                       
                            (tmr_registers(0)(70) and tmr_registers(2)(70));                                                         
                                                                                                                                     
        global_tmr_voter(1)(71)  <=    (tmr_registers(0)(71) and tmr_registers(1)(71)) or                                            
                            (tmr_registers(1)(71) and tmr_registers(2)(71)) or                                                       
                            (tmr_registers(0)(71) and tmr_registers(2)(71));                                                         
                                                                                                                                     
        global_tmr_voter(1)(72)  <=    (tmr_registers(0)(72) and tmr_registers(1)(72)) or                                            
                            (tmr_registers(1)(72) and tmr_registers(2)(72)) or                                                       
                            (tmr_registers(0)(72) and tmr_registers(2)(72));                                                         
                                                                                                                                     
        global_tmr_voter(1)(73)  <=    (tmr_registers(0)(73) and tmr_registers(1)(73)) or                                            
                            (tmr_registers(1)(73) and tmr_registers(2)(73)) or                                                       
                            (tmr_registers(0)(73) and tmr_registers(2)(73));                                                         
                                                                                                                                     
        global_tmr_voter(1)(74)  <=    (tmr_registers(0)(74) and tmr_registers(1)(74)) or                                            
                            (tmr_registers(1)(74) and tmr_registers(2)(74)) or                                                       
                            (tmr_registers(0)(74) and tmr_registers(2)(74));                                                         
                                                                                                                                     
        global_tmr_voter(1)(75)  <=    (tmr_registers(0)(75) and tmr_registers(1)(75)) or                                            
                            (tmr_registers(1)(75) and tmr_registers(2)(75)) or                                                       
                            (tmr_registers(0)(75) and tmr_registers(2)(75));                                                         
                                                                                                                                     
        global_tmr_voter(1)(76)  <=    (tmr_registers(0)(76) and tmr_registers(1)(76)) or                                            
                            (tmr_registers(1)(76) and tmr_registers(2)(76)) or                                                       
                            (tmr_registers(0)(76) and tmr_registers(2)(76));                                                         
                                                                                                                                     
        global_tmr_voter(1)(77)  <=    (tmr_registers(0)(77) and tmr_registers(1)(77)) or                                            
                            (tmr_registers(1)(77) and tmr_registers(2)(77)) or                                                       
                            (tmr_registers(0)(77) and tmr_registers(2)(77));                                                         
                                                                                                                                     
        global_tmr_voter(1)(78)  <=    (tmr_registers(0)(78) and tmr_registers(1)(78)) or                                            
                            (tmr_registers(1)(78) and tmr_registers(2)(78)) or                                                       
                            (tmr_registers(0)(78) and tmr_registers(2)(78));                                                         
                                                                                                                                     
        global_tmr_voter(1)(79)  <=    (tmr_registers(0)(79) and tmr_registers(1)(79)) or                                            
                            (tmr_registers(1)(79) and tmr_registers(2)(79)) or                                                       
                            (tmr_registers(0)(79) and tmr_registers(2)(79));                                                         
                                                                                                                                     
        global_tmr_voter(1)(80)  <=    (tmr_registers(0)(80) and tmr_registers(1)(80)) or                                            
                            (tmr_registers(1)(80) and tmr_registers(2)(80)) or                                                       
                            (tmr_registers(0)(80) and tmr_registers(2)(80));                                                         
                                                                                                                                     
        global_tmr_voter(1)(81)  <=    (tmr_registers(0)(81) and tmr_registers(1)(81)) or                                            
                            (tmr_registers(1)(81) and tmr_registers(2)(81)) or                                                       
                            (tmr_registers(0)(81) and tmr_registers(2)(81));                                                         
                                                                                                                                     
        global_tmr_voter(1)(82)  <=    (tmr_registers(0)(82) and tmr_registers(1)(82)) or                                            
                            (tmr_registers(1)(82) and tmr_registers(2)(82)) or                                                       
                            (tmr_registers(0)(82) and tmr_registers(2)(82));                                                         
                                                                                                                                     
        global_tmr_voter(1)(83)  <=    (tmr_registers(0)(83) and tmr_registers(1)(83)) or                                            
                            (tmr_registers(1)(83) and tmr_registers(2)(83)) or                                                       
                            (tmr_registers(0)(83) and tmr_registers(2)(83));                                                         
                                                                                                                                     
        global_tmr_voter(1)(84)  <=    (tmr_registers(0)(84) and tmr_registers(1)(84)) or                                            
                            (tmr_registers(1)(84) and tmr_registers(2)(84)) or                                                       
                            (tmr_registers(0)(84) and tmr_registers(2)(84));                                                         
                                                                                                                                     
        global_tmr_voter(1)(85)  <=    (tmr_registers(0)(85) and tmr_registers(1)(85)) or                                            
                            (tmr_registers(1)(85) and tmr_registers(2)(85)) or                                                       
                            (tmr_registers(0)(85) and tmr_registers(2)(85));                                                         
                                                                                                                                     
        global_tmr_voter(1)(86)  <=    (tmr_registers(0)(86) and tmr_registers(1)(86)) or                                            
                            (tmr_registers(1)(86) and tmr_registers(2)(86)) or                                                       
                            (tmr_registers(0)(86) and tmr_registers(2)(86));                                                         
                                                                                                                                     
        global_tmr_voter(1)(87)  <=    (tmr_registers(0)(87) and tmr_registers(1)(87)) or                                            
                            (tmr_registers(1)(87) and tmr_registers(2)(87)) or                                                       
                            (tmr_registers(0)(87) and tmr_registers(2)(87));                                                         
                                                                                                                                     
        global_tmr_voter(1)(88)  <=    (tmr_registers(0)(88) and tmr_registers(1)(88)) or                                            
                            (tmr_registers(1)(88) and tmr_registers(2)(88)) or                                                       
                            (tmr_registers(0)(88) and tmr_registers(2)(88));                                                         
                                                                                                                                     
        global_tmr_voter(1)(89)  <=    (tmr_registers(0)(89) and tmr_registers(1)(89)) or                                            
                            (tmr_registers(1)(89) and tmr_registers(2)(89)) or                                                       
                            (tmr_registers(0)(89) and tmr_registers(2)(89));                                                         
                                                                                                                                     
        global_tmr_voter(1)(90)  <=    (tmr_registers(0)(90) and tmr_registers(1)(90)) or                                            
                            (tmr_registers(1)(90) and tmr_registers(2)(90)) or                                                       
                            (tmr_registers(0)(90) and tmr_registers(2)(90));                                                         
                                                                                                                                     
        global_tmr_voter(1)(91)  <=    (tmr_registers(0)(91) and tmr_registers(1)(91)) or                                            
                            (tmr_registers(1)(91) and tmr_registers(2)(91)) or                                                       
                            (tmr_registers(0)(91) and tmr_registers(2)(91));                                                         
                                                                                                                                     
        global_tmr_voter(1)(92)  <=    (tmr_registers(0)(92) and tmr_registers(1)(92)) or                                            
                            (tmr_registers(1)(92) and tmr_registers(2)(92)) or                                                       
                            (tmr_registers(0)(92) and tmr_registers(2)(92));                                                         
                                                                                                                                     
        global_tmr_voter(1)(93)  <=    (tmr_registers(0)(93) and tmr_registers(1)(93)) or                                            
                            (tmr_registers(1)(93) and tmr_registers(2)(93)) or                                                       
                            (tmr_registers(0)(93) and tmr_registers(2)(93));                                                         
                                                                                                                                     
        global_tmr_voter(1)(94)  <=    (tmr_registers(0)(94) and tmr_registers(1)(94)) or                                            
                            (tmr_registers(1)(94) and tmr_registers(2)(94)) or                                                       
                            (tmr_registers(0)(94) and tmr_registers(2)(94));                                                         
                                                                                                                                     
        global_tmr_voter(1)(95)  <=    (tmr_registers(0)(95) and tmr_registers(1)(95)) or                                            
                            (tmr_registers(1)(95) and tmr_registers(2)(95)) or                                                       
                            (tmr_registers(0)(95) and tmr_registers(2)(95));                                                         
                                                                                                                                     
        global_tmr_voter(1)(96)  <=    (tmr_registers(0)(96) and tmr_registers(1)(96)) or                                            
                            (tmr_registers(1)(96) and tmr_registers(2)(96)) or                                                       
                            (tmr_registers(0)(96) and tmr_registers(2)(96));                                                         
                                                                                                                                     
        global_tmr_voter(1)(97)  <=    (tmr_registers(0)(97) and tmr_registers(1)(97)) or                                            
                            (tmr_registers(1)(97) and tmr_registers(2)(97)) or                                                       
                            (tmr_registers(0)(97) and tmr_registers(2)(97));                                                         
                                                                                                                                     
        global_tmr_voter(1)(98)  <=    (tmr_registers(0)(98) and tmr_registers(1)(98)) or                                            
                            (tmr_registers(1)(98) and tmr_registers(2)(98)) or                                                       
                            (tmr_registers(0)(98) and tmr_registers(2)(98));                                                         
                                                                                                                                     
        global_tmr_voter(1)(99)  <=    (tmr_registers(0)(99) and tmr_registers(1)(99)) or                                            
                            (tmr_registers(1)(99) and tmr_registers(2)(99)) or                                                       
                            (tmr_registers(0)(99) and tmr_registers(2)(99));                                                         
                                                                                                                                     
        global_tmr_voter(1)(100)  <=    (tmr_registers(0)(100) and tmr_registers(1)(100)) or                                            
                            (tmr_registers(1)(100) and tmr_registers(2)(100)) or                                                       
                            (tmr_registers(0)(100) and tmr_registers(2)(100));                                                         
                                                                                                                                     
        global_tmr_voter(1)(101)  <=    (tmr_registers(0)(101) and tmr_registers(1)(101)) or                                            
                            (tmr_registers(1)(101) and tmr_registers(2)(101)) or                                                       
                            (tmr_registers(0)(101) and tmr_registers(2)(101));                                                         
                                                                                                                                     
        global_tmr_voter(1)(102)  <=    (tmr_registers(0)(102) and tmr_registers(1)(102)) or                                            
                            (tmr_registers(1)(102) and tmr_registers(2)(102)) or                                                       
                            (tmr_registers(0)(102) and tmr_registers(2)(102));                                                         
                                                                                                                                     
        global_tmr_voter(1)(103)  <=    (tmr_registers(0)(103) and tmr_registers(1)(103)) or                                            
                            (tmr_registers(1)(103) and tmr_registers(2)(103)) or                                                       
                            (tmr_registers(0)(103) and tmr_registers(2)(103));                                                         
                                                                                                                                     
        global_tmr_voter(1)(104)  <=    (tmr_registers(0)(104) and tmr_registers(1)(104)) or                                            
                            (tmr_registers(1)(104) and tmr_registers(2)(104)) or                                                       
                            (tmr_registers(0)(104) and tmr_registers(2)(104));                                                         
                                                                                                                                     
        global_tmr_voter(1)(105)  <=    (tmr_registers(0)(105) and tmr_registers(1)(105)) or                                            
                            (tmr_registers(1)(105) and tmr_registers(2)(105)) or                                                       
                            (tmr_registers(0)(105) and tmr_registers(2)(105));                                                         
                                                                                                                                     
        global_tmr_voter(1)(106)  <=    (tmr_registers(0)(106) and tmr_registers(1)(106)) or                                            
                            (tmr_registers(1)(106) and tmr_registers(2)(106)) or                                                       
                            (tmr_registers(0)(106) and tmr_registers(2)(106));                                                         
                                                                                                                                     
        global_tmr_voter(1)(107)  <=    (tmr_registers(0)(107) and tmr_registers(1)(107)) or                                            
                            (tmr_registers(1)(107) and tmr_registers(2)(107)) or                                                       
                            (tmr_registers(0)(107) and tmr_registers(2)(107));                                                         
                                                                                                                                     
        global_tmr_voter(1)(108)  <=    (tmr_registers(0)(108) and tmr_registers(1)(108)) or                                            
                            (tmr_registers(1)(108) and tmr_registers(2)(108)) or                                                       
                            (tmr_registers(0)(108) and tmr_registers(2)(108));                                                         
                                                                                                                                     
        global_tmr_voter(1)(109)  <=    (tmr_registers(0)(109) and tmr_registers(1)(109)) or                                            
                            (tmr_registers(1)(109) and tmr_registers(2)(109)) or                                                       
                            (tmr_registers(0)(109) and tmr_registers(2)(109));                                                         
                                                                                                                                     
        global_tmr_voter(1)(110)  <=    (tmr_registers(0)(110) and tmr_registers(1)(110)) or                                            
                            (tmr_registers(1)(110) and tmr_registers(2)(110)) or                                                       
                            (tmr_registers(0)(110) and tmr_registers(2)(110));                                                         
                                                                                                                                     
        global_tmr_voter(1)(111)  <=    (tmr_registers(0)(111) and tmr_registers(1)(111)) or                                            
                            (tmr_registers(1)(111) and tmr_registers(2)(111)) or                                                       
                            (tmr_registers(0)(111) and tmr_registers(2)(111));                                                         
                                                                                                                                     
        global_tmr_voter(1)(112)  <=    (tmr_registers(0)(112) and tmr_registers(1)(112)) or                                            
                            (tmr_registers(1)(112) and tmr_registers(2)(112)) or                                                       
                            (tmr_registers(0)(112) and tmr_registers(2)(112));                                                         
                                                                                                                                     
        global_tmr_voter(1)(113)  <=    (tmr_registers(0)(113) and tmr_registers(1)(113)) or                                            
                            (tmr_registers(1)(113) and tmr_registers(2)(113)) or                                                       
                            (tmr_registers(0)(113) and tmr_registers(2)(113));                                                         
                                                                                                                                     
        global_tmr_voter(1)(114)  <=    (tmr_registers(0)(114) and tmr_registers(1)(114)) or                                            
                            (tmr_registers(1)(114) and tmr_registers(2)(114)) or                                                       
                            (tmr_registers(0)(114) and tmr_registers(2)(114));                                                         
                                                                                                                                     
        global_tmr_voter(1)(115)  <=    (tmr_registers(0)(115) and tmr_registers(1)(115)) or                                            
                            (tmr_registers(1)(115) and tmr_registers(2)(115)) or                                                       
                            (tmr_registers(0)(115) and tmr_registers(2)(115));                                                         
                                                                                                                                     
        global_tmr_voter(1)(116)  <=    (tmr_registers(0)(116) and tmr_registers(1)(116)) or                                            
                            (tmr_registers(1)(116) and tmr_registers(2)(116)) or                                                       
                            (tmr_registers(0)(116) and tmr_registers(2)(116));                                                         
                                                                                                                                     
        global_tmr_voter(1)(117)  <=    (tmr_registers(0)(117) and tmr_registers(1)(117)) or                                            
                            (tmr_registers(1)(117) and tmr_registers(2)(117)) or                                                       
                            (tmr_registers(0)(117) and tmr_registers(2)(117));                                                         
                                                                                                                                     
        global_tmr_voter(1)(118)  <=    (tmr_registers(0)(118) and tmr_registers(1)(118)) or                                            
                            (tmr_registers(1)(118) and tmr_registers(2)(118)) or                                                       
                            (tmr_registers(0)(118) and tmr_registers(2)(118));                                                         
                                                                                                                                     
        global_tmr_voter(1)(119)  <=    (tmr_registers(0)(119) and tmr_registers(1)(119)) or                                            
                            (tmr_registers(1)(119) and tmr_registers(2)(119)) or                                                       
                            (tmr_registers(0)(119) and tmr_registers(2)(119));                                                         
                                                                                                                                     
        global_tmr_voter(1)(120)  <=    (tmr_registers(0)(120) and tmr_registers(1)(120)) or                                            
                            (tmr_registers(1)(120) and tmr_registers(2)(120)) or                                                       
                            (tmr_registers(0)(120) and tmr_registers(2)(120));                                                         
                                                                                                                                     
        global_tmr_voter(1)(121)  <=    (tmr_registers(0)(121) and tmr_registers(1)(121)) or                                            
                            (tmr_registers(1)(121) and tmr_registers(2)(121)) or                                                       
                            (tmr_registers(0)(121) and tmr_registers(2)(121));                                                         
                                                                                                                                     
        global_tmr_voter(1)(122)  <=    (tmr_registers(0)(122) and tmr_registers(1)(122)) or                                            
                            (tmr_registers(1)(122) and tmr_registers(2)(122)) or                                                       
                            (tmr_registers(0)(122) and tmr_registers(2)(122));                                                         
                                                                                                                                     
        global_tmr_voter(1)(123)  <=    (tmr_registers(0)(123) and tmr_registers(1)(123)) or                                            
                            (tmr_registers(1)(123) and tmr_registers(2)(123)) or                                                       
                            (tmr_registers(0)(123) and tmr_registers(2)(123));                                                         
                                                                                                                                     
        global_tmr_voter(1)(124)  <=    (tmr_registers(0)(124) and tmr_registers(1)(124)) or                                            
                            (tmr_registers(1)(124) and tmr_registers(2)(124)) or                                                       
                            (tmr_registers(0)(124) and tmr_registers(2)(124));                                                         
                                                                                                                                     
        global_tmr_voter(1)(125)  <=    (tmr_registers(0)(125) and tmr_registers(1)(125)) or                                            
                            (tmr_registers(1)(125) and tmr_registers(2)(125)) or                                                       
                            (tmr_registers(0)(125) and tmr_registers(2)(125));                                                         
                                                                                                                                     
        global_tmr_voter(1)(126)  <=    (tmr_registers(0)(126) and tmr_registers(1)(126)) or                                            
                            (tmr_registers(1)(126) and tmr_registers(2)(126)) or                                                       
                            (tmr_registers(0)(126) and tmr_registers(2)(126));                                                         
                                                                                                                                     
        global_tmr_voter(1)(127)  <=    (tmr_registers(0)(127) and tmr_registers(1)(127)) or                                            
                            (tmr_registers(1)(127) and tmr_registers(2)(127)) or                                                       
                            (tmr_registers(0)(127) and tmr_registers(2)(127));                                                         
                                                                                                                                     
        global_tmr_voter(1)(128)  <=    (tmr_registers(0)(128) and tmr_registers(1)(128)) or                                            
                            (tmr_registers(1)(128) and tmr_registers(2)(128)) or                                                       
                            (tmr_registers(0)(128) and tmr_registers(2)(128));                                                         
                                                                                                                                     
        global_tmr_voter(1)(129)  <=    (tmr_registers(0)(129) and tmr_registers(1)(129)) or                                            
                            (tmr_registers(1)(129) and tmr_registers(2)(129)) or                                                       
                            (tmr_registers(0)(129) and tmr_registers(2)(129));                                                         
                                                                                                                                     
        global_tmr_voter(1)(130)  <=    (tmr_registers(0)(130) and tmr_registers(1)(130)) or                                            
                            (tmr_registers(1)(130) and tmr_registers(2)(130)) or                                                       
                            (tmr_registers(0)(130) and tmr_registers(2)(130));                                                         
                                                                                                                                     
        global_tmr_voter(1)(131)  <=    (tmr_registers(0)(131) and tmr_registers(1)(131)) or                                            
                            (tmr_registers(1)(131) and tmr_registers(2)(131)) or                                                       
                            (tmr_registers(0)(131) and tmr_registers(2)(131));                                                         
                                                                                                                                     
        global_tmr_voter(1)(132)  <=    (tmr_registers(0)(132) and tmr_registers(1)(132)) or                                            
                            (tmr_registers(1)(132) and tmr_registers(2)(132)) or                                                       
                            (tmr_registers(0)(132) and tmr_registers(2)(132));                                                         
                                                                                                                                     
        global_tmr_voter(1)(133)  <=    (tmr_registers(0)(133) and tmr_registers(1)(133)) or                                            
                            (tmr_registers(1)(133) and tmr_registers(2)(133)) or                                                       
                            (tmr_registers(0)(133) and tmr_registers(2)(133));                                                         
                                                                                                                                     
        global_tmr_voter(1)(134)  <=    (tmr_registers(0)(134) and tmr_registers(1)(134)) or                                            
                            (tmr_registers(1)(134) and tmr_registers(2)(134)) or                                                       
                            (tmr_registers(0)(134) and tmr_registers(2)(134));                                                         
                                                                                                                                     
        global_tmr_voter(1)(135)  <=    (tmr_registers(0)(135) and tmr_registers(1)(135)) or                                            
                            (tmr_registers(1)(135) and tmr_registers(2)(135)) or                                                       
                            (tmr_registers(0)(135) and tmr_registers(2)(135));                                                         
                                                                                                                                     
        global_tmr_voter(1)(136)  <=    (tmr_registers(0)(136) and tmr_registers(1)(136)) or                                            
                            (tmr_registers(1)(136) and tmr_registers(2)(136)) or                                                       
                            (tmr_registers(0)(136) and tmr_registers(2)(136));                                                         
                                                                                                                                     
        global_tmr_voter(1)(137)  <=    (tmr_registers(0)(137) and tmr_registers(1)(137)) or                                            
                            (tmr_registers(1)(137) and tmr_registers(2)(137)) or                                                       
                            (tmr_registers(0)(137) and tmr_registers(2)(137));                                                         
                                                                                                                                     
        global_tmr_voter(1)(138)  <=    (tmr_registers(0)(138) and tmr_registers(1)(138)) or                                            
                            (tmr_registers(1)(138) and tmr_registers(2)(138)) or                                                       
                            (tmr_registers(0)(138) and tmr_registers(2)(138));                                                         
                                                                                                                                     
        global_tmr_voter(1)(139)  <=    (tmr_registers(0)(139) and tmr_registers(1)(139)) or                                            
                            (tmr_registers(1)(139) and tmr_registers(2)(139)) or                                                       
                            (tmr_registers(0)(139) and tmr_registers(2)(139));                                                         
                                                                                                                                     
        global_tmr_voter(1)(140)  <=    (tmr_registers(0)(140) and tmr_registers(1)(140)) or                                            
                            (tmr_registers(1)(140) and tmr_registers(2)(140)) or                                                       
                            (tmr_registers(0)(140) and tmr_registers(2)(140));                                                         
                                                                                                                                     
        global_tmr_voter(1)(141)  <=    (tmr_registers(0)(141) and tmr_registers(1)(141)) or                                            
                            (tmr_registers(1)(141) and tmr_registers(2)(141)) or                                                       
                            (tmr_registers(0)(141) and tmr_registers(2)(141));                                                         
                                                                                                                                     
        global_tmr_voter(1)(142)  <=    (tmr_registers(0)(142) and tmr_registers(1)(142)) or                                            
                            (tmr_registers(1)(142) and tmr_registers(2)(142)) or                                                       
                            (tmr_registers(0)(142) and tmr_registers(2)(142));                                                         
                                                                                                                                     
        global_tmr_voter(1)(143)  <=    (tmr_registers(0)(143) and tmr_registers(1)(143)) or                                            
                            (tmr_registers(1)(143) and tmr_registers(2)(143)) or                                                       
                            (tmr_registers(0)(143) and tmr_registers(2)(143));                                                         
                                                                                                                                     
        global_tmr_voter(1)(144)  <=    (tmr_registers(0)(144) and tmr_registers(1)(144)) or                                            
                            (tmr_registers(1)(144) and tmr_registers(2)(144)) or                                                       
                            (tmr_registers(0)(144) and tmr_registers(2)(144));                                                         
                                                                                                                                     
        global_tmr_voter(1)(145)  <=    (tmr_registers(0)(145) and tmr_registers(1)(145)) or                                            
                            (tmr_registers(1)(145) and tmr_registers(2)(145)) or                                                       
                            (tmr_registers(0)(145) and tmr_registers(2)(145));                                                         
                                                                                                                                     
        global_tmr_voter(1)(146)  <=    (tmr_registers(0)(146) and tmr_registers(1)(146)) or                                            
                            (tmr_registers(1)(146) and tmr_registers(2)(146)) or                                                       
                            (tmr_registers(0)(146) and tmr_registers(2)(146));                                                         
                                                                                                                                     
        global_tmr_voter(1)(147)  <=    (tmr_registers(0)(147) and tmr_registers(1)(147)) or                                            
                            (tmr_registers(1)(147) and tmr_registers(2)(147)) or                                                       
                            (tmr_registers(0)(147) and tmr_registers(2)(147));                                                         
                                                                                                                                     
        global_tmr_voter(1)(148)  <=    (tmr_registers(0)(148) and tmr_registers(1)(148)) or                                            
                            (tmr_registers(1)(148) and tmr_registers(2)(148)) or                                                       
                            (tmr_registers(0)(148) and tmr_registers(2)(148));                                                         
                                                                                                                                     
        global_tmr_voter(1)(149)  <=    (tmr_registers(0)(149) and tmr_registers(1)(149)) or                                            
                            (tmr_registers(1)(149) and tmr_registers(2)(149)) or                                                       
                            (tmr_registers(0)(149) and tmr_registers(2)(149));                                                         
                                                                                                                                     
        global_tmr_voter(1)(150)  <=    (tmr_registers(0)(150) and tmr_registers(1)(150)) or                                            
                            (tmr_registers(1)(150) and tmr_registers(2)(150)) or                                                       
                            (tmr_registers(0)(150) and tmr_registers(2)(150));                                                         
                                                                                                                                     
        global_tmr_voter(1)(151)  <=    (tmr_registers(0)(151) and tmr_registers(1)(151)) or                                            
                            (tmr_registers(1)(151) and tmr_registers(2)(151)) or                                                       
                            (tmr_registers(0)(151) and tmr_registers(2)(151));                                                         
                                                                                                                                     
        global_tmr_voter(1)(152)  <=    (tmr_registers(0)(152) and tmr_registers(1)(152)) or                                            
                            (tmr_registers(1)(152) and tmr_registers(2)(152)) or                                                       
                            (tmr_registers(0)(152) and tmr_registers(2)(152));                                                         
                                                                                                                                     
        global_tmr_voter(1)(153)  <=    (tmr_registers(0)(153) and tmr_registers(1)(153)) or                                            
                            (tmr_registers(1)(153) and tmr_registers(2)(153)) or                                                       
                            (tmr_registers(0)(153) and tmr_registers(2)(153));                                                         
                                                                                                                                     
        global_tmr_voter(1)(154)  <=    (tmr_registers(0)(154) and tmr_registers(1)(154)) or                                            
                            (tmr_registers(1)(154) and tmr_registers(2)(154)) or                                                       
                            (tmr_registers(0)(154) and tmr_registers(2)(154));                                                         
                                                                                                                                     
        global_tmr_voter(1)(155)  <=    (tmr_registers(0)(155) and tmr_registers(1)(155)) or                                            
                            (tmr_registers(1)(155) and tmr_registers(2)(155)) or                                                       
                            (tmr_registers(0)(155) and tmr_registers(2)(155));                                                         
                                                                                                                                     
        global_tmr_voter(1)(156)  <=    (tmr_registers(0)(156) and tmr_registers(1)(156)) or                                            
                            (tmr_registers(1)(156) and tmr_registers(2)(156)) or                                                       
                            (tmr_registers(0)(156) and tmr_registers(2)(156));                                                         
                                                                                                                                     
        global_tmr_voter(1)(157)  <=    (tmr_registers(0)(157) and tmr_registers(1)(157)) or                                            
                            (tmr_registers(1)(157) and tmr_registers(2)(157)) or                                                       
                            (tmr_registers(0)(157) and tmr_registers(2)(157));                                                         
                                                                                                                                     
        global_tmr_voter(1)(158)  <=    (tmr_registers(0)(158) and tmr_registers(1)(158)) or                                            
                            (tmr_registers(1)(158) and tmr_registers(2)(158)) or                                                       
                            (tmr_registers(0)(158) and tmr_registers(2)(158));                                                         
                                                                                                                                     
        global_tmr_voter(1)(159)  <=    (tmr_registers(0)(159) and tmr_registers(1)(159)) or                                            
                            (tmr_registers(1)(159) and tmr_registers(2)(159)) or                                                       
                            (tmr_registers(0)(159) and tmr_registers(2)(159));                                                         
                                                                                                                                     
        global_tmr_voter(1)(160)  <=    (tmr_registers(0)(160) and tmr_registers(1)(160)) or                                            
                            (tmr_registers(1)(160) and tmr_registers(2)(160)) or                                                       
                            (tmr_registers(0)(160) and tmr_registers(2)(160));                                                         
                                                                                                                                     
        global_tmr_voter(1)(161)  <=    (tmr_registers(0)(161) and tmr_registers(1)(161)) or                                            
                            (tmr_registers(1)(161) and tmr_registers(2)(161)) or                                                       
                            (tmr_registers(0)(161) and tmr_registers(2)(161));                                                         
                                                                                                                                     
        global_tmr_voter(1)(162)  <=    (tmr_registers(0)(162) and tmr_registers(1)(162)) or                                            
                            (tmr_registers(1)(162) and tmr_registers(2)(162)) or                                                       
                            (tmr_registers(0)(162) and tmr_registers(2)(162));                                                         
                                                                                                                                     
        global_tmr_voter(1)(163)  <=    (tmr_registers(0)(163) and tmr_registers(1)(163)) or                                            
                            (tmr_registers(1)(163) and tmr_registers(2)(163)) or                                                       
                            (tmr_registers(0)(163) and tmr_registers(2)(163));                                                         
                                                                                                                                     
        global_tmr_voter(1)(164)  <=    (tmr_registers(0)(164) and tmr_registers(1)(164)) or                                            
                            (tmr_registers(1)(164) and tmr_registers(2)(164)) or                                                       
                            (tmr_registers(0)(164) and tmr_registers(2)(164));                                                         
                                                                                                                                     
        global_tmr_voter(1)(165)  <=    (tmr_registers(0)(165) and tmr_registers(1)(165)) or                                            
                            (tmr_registers(1)(165) and tmr_registers(2)(165)) or                                                       
                            (tmr_registers(0)(165) and tmr_registers(2)(165));                                                         
                                                                                                                                     
        global_tmr_voter(1)(166)  <=    (tmr_registers(0)(166) and tmr_registers(1)(166)) or                                            
                            (tmr_registers(1)(166) and tmr_registers(2)(166)) or                                                       
                            (tmr_registers(0)(166) and tmr_registers(2)(166));                                                         
                                                                                                                                     
        global_tmr_voter(1)(167)  <=    (tmr_registers(0)(167) and tmr_registers(1)(167)) or                                            
                            (tmr_registers(1)(167) and tmr_registers(2)(167)) or                                                       
                            (tmr_registers(0)(167) and tmr_registers(2)(167));                                                         
                                                                                                                                     
        global_tmr_voter(1)(168)  <=    (tmr_registers(0)(168) and tmr_registers(1)(168)) or                                            
                            (tmr_registers(1)(168) and tmr_registers(2)(168)) or                                                       
                            (tmr_registers(0)(168) and tmr_registers(2)(168));                                                         
                                                                                                                                     
        global_tmr_voter(1)(169)  <=    (tmr_registers(0)(169) and tmr_registers(1)(169)) or                                            
                            (tmr_registers(1)(169) and tmr_registers(2)(169)) or                                                       
                            (tmr_registers(0)(169) and tmr_registers(2)(169));                                                         
                                                                                                                                     
        global_tmr_voter(1)(170)  <=    (tmr_registers(0)(170) and tmr_registers(1)(170)) or                                            
                            (tmr_registers(1)(170) and tmr_registers(2)(170)) or                                                       
                            (tmr_registers(0)(170) and tmr_registers(2)(170));                                                         
                                                                                                                                     
        global_tmr_voter(1)(171)  <=    (tmr_registers(0)(171) and tmr_registers(1)(171)) or                                            
                            (tmr_registers(1)(171) and tmr_registers(2)(171)) or                                                       
                            (tmr_registers(0)(171) and tmr_registers(2)(171));                                                         
                                                                                                                                     
        global_tmr_voter(1)(172)  <=    (tmr_registers(0)(172) and tmr_registers(1)(172)) or                                            
                            (tmr_registers(1)(172) and tmr_registers(2)(172)) or                                                       
                            (tmr_registers(0)(172) and tmr_registers(2)(172));                                                         
                                                                                                                                     
        global_tmr_voter(1)(173)  <=    (tmr_registers(0)(173) and tmr_registers(1)(173)) or                                            
                            (tmr_registers(1)(173) and tmr_registers(2)(173)) or                                                       
                            (tmr_registers(0)(173) and tmr_registers(2)(173));                                                         
                                                                                                                                     
        global_tmr_voter(1)(174)  <=    (tmr_registers(0)(174) and tmr_registers(1)(174)) or                                            
                            (tmr_registers(1)(174) and tmr_registers(2)(174)) or                                                       
                            (tmr_registers(0)(174) and tmr_registers(2)(174));                                                         
                                                                                                                                     
        global_tmr_voter(1)(175)  <=    (tmr_registers(0)(175) and tmr_registers(1)(175)) or                                            
                            (tmr_registers(1)(175) and tmr_registers(2)(175)) or                                                       
                            (tmr_registers(0)(175) and tmr_registers(2)(175));                                                         
                                                                                                                                     
        global_tmr_voter(1)(176)  <=    (tmr_registers(0)(176) and tmr_registers(1)(176)) or                                            
                            (tmr_registers(1)(176) and tmr_registers(2)(176)) or                                                       
                            (tmr_registers(0)(176) and tmr_registers(2)(176));                                                         
                                                                                                                                     
        global_tmr_voter(1)(177)  <=    (tmr_registers(0)(177) and tmr_registers(1)(177)) or                                            
                            (tmr_registers(1)(177) and tmr_registers(2)(177)) or                                                       
                            (tmr_registers(0)(177) and tmr_registers(2)(177));                                                         
                                                                                                                                     
        global_tmr_voter(1)(178)  <=    (tmr_registers(0)(178) and tmr_registers(1)(178)) or                                            
                            (tmr_registers(1)(178) and tmr_registers(2)(178)) or                                                       
                            (tmr_registers(0)(178) and tmr_registers(2)(178));                                                         
                                                                                                                                     
        global_tmr_voter(1)(179)  <=    (tmr_registers(0)(179) and tmr_registers(1)(179)) or                                            
                            (tmr_registers(1)(179) and tmr_registers(2)(179)) or                                                       
                            (tmr_registers(0)(179) and tmr_registers(2)(179));                                                         
                                                                                                                                     
        global_tmr_voter(1)(180)  <=    (tmr_registers(0)(180) and tmr_registers(1)(180)) or                                            
                            (tmr_registers(1)(180) and tmr_registers(2)(180)) or                                                       
                            (tmr_registers(0)(180) and tmr_registers(2)(180));                                                         
                                                                                                                                     
        global_tmr_voter(1)(181)  <=    (tmr_registers(0)(181) and tmr_registers(1)(181)) or                                            
                            (tmr_registers(1)(181) and tmr_registers(2)(181)) or                                                       
                            (tmr_registers(0)(181) and tmr_registers(2)(181));                                                         
                                                                                                                                     
        global_tmr_voter(1)(182)  <=    (tmr_registers(0)(182) and tmr_registers(1)(182)) or                                            
                            (tmr_registers(1)(182) and tmr_registers(2)(182)) or                                                       
                            (tmr_registers(0)(182) and tmr_registers(2)(182));                                                         
                                                                                                                                     
        global_tmr_voter(1)(183)  <=    (tmr_registers(0)(183) and tmr_registers(1)(183)) or                                            
                            (tmr_registers(1)(183) and tmr_registers(2)(183)) or                                                       
                            (tmr_registers(0)(183) and tmr_registers(2)(183));                                                         
                                                                                                                                     
        global_tmr_voter(1)(184)  <=    (tmr_registers(0)(184) and tmr_registers(1)(184)) or                                            
                            (tmr_registers(1)(184) and tmr_registers(2)(184)) or                                                       
                            (tmr_registers(0)(184) and tmr_registers(2)(184));                                                         
                                                                                                                                     
        global_tmr_voter(1)(185)  <=    (tmr_registers(0)(185) and tmr_registers(1)(185)) or                                            
                            (tmr_registers(1)(185) and tmr_registers(2)(185)) or                                                       
                            (tmr_registers(0)(185) and tmr_registers(2)(185));                                                         
                                                                                                                                     
        global_tmr_voter(1)(186)  <=    (tmr_registers(0)(186) and tmr_registers(1)(186)) or                                            
                            (tmr_registers(1)(186) and tmr_registers(2)(186)) or                                                       
                            (tmr_registers(0)(186) and tmr_registers(2)(186));                                                         
                                                                                                                                     
        global_tmr_voter(1)(187)  <=    (tmr_registers(0)(187) and tmr_registers(1)(187)) or                                            
                            (tmr_registers(1)(187) and tmr_registers(2)(187)) or                                                       
                            (tmr_registers(0)(187) and tmr_registers(2)(187));                                                         
                                                                                                                                     
        global_tmr_voter(1)(188)  <=    (tmr_registers(0)(188) and tmr_registers(1)(188)) or                                            
                            (tmr_registers(1)(188) and tmr_registers(2)(188)) or                                                       
                            (tmr_registers(0)(188) and tmr_registers(2)(188));                                                         
                                                                                                                                     
        global_tmr_voter(1)(189)  <=    (tmr_registers(0)(189) and tmr_registers(1)(189)) or                                            
                            (tmr_registers(1)(189) and tmr_registers(2)(189)) or                                                       
                            (tmr_registers(0)(189) and tmr_registers(2)(189));                                                         
                                                                                                                                     
        global_tmr_voter(1)(190)  <=    (tmr_registers(0)(190) and tmr_registers(1)(190)) or                                            
                            (tmr_registers(1)(190) and tmr_registers(2)(190)) or                                                       
                            (tmr_registers(0)(190) and tmr_registers(2)(190));                                                         
                                                                                                                                     
        global_tmr_voter(1)(191)  <=    (tmr_registers(0)(191) and tmr_registers(1)(191)) or                                            
                            (tmr_registers(1)(191) and tmr_registers(2)(191)) or                                                       
                            (tmr_registers(0)(191) and tmr_registers(2)(191));                                                         
                                                                                                                                     
        global_tmr_voter(1)(192)  <=    (tmr_registers(0)(192) and tmr_registers(1)(192)) or                                            
                            (tmr_registers(1)(192) and tmr_registers(2)(192)) or                                                       
                            (tmr_registers(0)(192) and tmr_registers(2)(192));                                                         
                                                                                                                                     
        global_tmr_voter(1)(193)  <=    (tmr_registers(0)(193) and tmr_registers(1)(193)) or                                            
                            (tmr_registers(1)(193) and tmr_registers(2)(193)) or                                                       
                            (tmr_registers(0)(193) and tmr_registers(2)(193));                                                         
                                                                                                                                     
        global_tmr_voter(1)(194)  <=    (tmr_registers(0)(194) and tmr_registers(1)(194)) or                                            
                            (tmr_registers(1)(194) and tmr_registers(2)(194)) or                                                       
                            (tmr_registers(0)(194) and tmr_registers(2)(194));                                                         
                                                                                                                                     
        global_tmr_voter(1)(195)  <=    (tmr_registers(0)(195) and tmr_registers(1)(195)) or                                            
                            (tmr_registers(1)(195) and tmr_registers(2)(195)) or                                                       
                            (tmr_registers(0)(195) and tmr_registers(2)(195));                                                         
                                                                                                                                     
        global_tmr_voter(1)(196)  <=    (tmr_registers(0)(196) and tmr_registers(1)(196)) or                                            
                            (tmr_registers(1)(196) and tmr_registers(2)(196)) or                                                       
                            (tmr_registers(0)(196) and tmr_registers(2)(196));                                                         
                                                                                                                                     
        global_tmr_voter(1)(197)  <=    (tmr_registers(0)(197) and tmr_registers(1)(197)) or                                            
                            (tmr_registers(1)(197) and tmr_registers(2)(197)) or                                                       
                            (tmr_registers(0)(197) and tmr_registers(2)(197));                                                         
                                                                                                                                     
        global_tmr_voter(1)(198)  <=    (tmr_registers(0)(198) and tmr_registers(1)(198)) or                                            
                            (tmr_registers(1)(198) and tmr_registers(2)(198)) or                                                       
                            (tmr_registers(0)(198) and tmr_registers(2)(198));                                                         
                                                                                                                                     
        global_tmr_voter(1)(199)  <=    (tmr_registers(0)(199) and tmr_registers(1)(199)) or                                            
                            (tmr_registers(1)(199) and tmr_registers(2)(199)) or                                                       
                            (tmr_registers(0)(199) and tmr_registers(2)(199));                                                         
                                                                                                                                     
        global_tmr_voter(1)(200)  <=    (tmr_registers(0)(200) and tmr_registers(1)(200)) or                                            
                            (tmr_registers(1)(200) and tmr_registers(2)(200)) or                                                       
                            (tmr_registers(0)(200) and tmr_registers(2)(200));                                                         
                                                                                                                                     
        global_tmr_voter(1)(201)  <=    (tmr_registers(0)(201) and tmr_registers(1)(201)) or                                            
                            (tmr_registers(1)(201) and tmr_registers(2)(201)) or                                                       
                            (tmr_registers(0)(201) and tmr_registers(2)(201));                                                         
                                                                                                                                     
        global_tmr_voter(1)(202)  <=    (tmr_registers(0)(202) and tmr_registers(1)(202)) or                                            
                            (tmr_registers(1)(202) and tmr_registers(2)(202)) or                                                       
                            (tmr_registers(0)(202) and tmr_registers(2)(202));                                                         
                                                                                                                                     
        global_tmr_voter(1)(203)  <=    (tmr_registers(0)(203) and tmr_registers(1)(203)) or                                            
                            (tmr_registers(1)(203) and tmr_registers(2)(203)) or                                                       
                            (tmr_registers(0)(203) and tmr_registers(2)(203));                                                         
                                                                                                                                     
        global_tmr_voter(1)(204)  <=    (tmr_registers(0)(204) and tmr_registers(1)(204)) or                                            
                            (tmr_registers(1)(204) and tmr_registers(2)(204)) or                                                       
                            (tmr_registers(0)(204) and tmr_registers(2)(204));                                                         
                                                                                                                                     
        global_tmr_voter(1)(205)  <=    (tmr_registers(0)(205) and tmr_registers(1)(205)) or                                            
                            (tmr_registers(1)(205) and tmr_registers(2)(205)) or                                                       
                            (tmr_registers(0)(205) and tmr_registers(2)(205));                                                         
                                                                                                                                     
        global_tmr_voter(1)(206)  <=    (tmr_registers(0)(206) and tmr_registers(1)(206)) or                                            
                            (tmr_registers(1)(206) and tmr_registers(2)(206)) or                                                       
                            (tmr_registers(0)(206) and tmr_registers(2)(206));                                                         
                                                                                                                                     
        global_tmr_voter(1)(207)  <=    (tmr_registers(0)(207) and tmr_registers(1)(207)) or                                            
                            (tmr_registers(1)(207) and tmr_registers(2)(207)) or                                                       
                            (tmr_registers(0)(207) and tmr_registers(2)(207));                                                         
                                                                                                                                     
        global_tmr_voter(1)(208)  <=    (tmr_registers(0)(208) and tmr_registers(1)(208)) or                                            
                            (tmr_registers(1)(208) and tmr_registers(2)(208)) or                                                       
                            (tmr_registers(0)(208) and tmr_registers(2)(208));                                                         
                                                                                                                                     
        global_tmr_voter(1)(209)  <=    (tmr_registers(0)(209) and tmr_registers(1)(209)) or                                            
                            (tmr_registers(1)(209) and tmr_registers(2)(209)) or                                                       
                            (tmr_registers(0)(209) and tmr_registers(2)(209));                                                         
                                                                                                                                     
        global_tmr_voter(1)(210)  <=    (tmr_registers(0)(210) and tmr_registers(1)(210)) or                                            
                            (tmr_registers(1)(210) and tmr_registers(2)(210)) or                                                       
                            (tmr_registers(0)(210) and tmr_registers(2)(210));                                                         
                                                                                                                                     
        global_tmr_voter(1)(211)  <=    (tmr_registers(0)(211) and tmr_registers(1)(211)) or                                            
                            (tmr_registers(1)(211) and tmr_registers(2)(211)) or                                                       
                            (tmr_registers(0)(211) and tmr_registers(2)(211));                                                         
                                                                                                                                     
        global_tmr_voter(1)(212)  <=    (tmr_registers(0)(212) and tmr_registers(1)(212)) or                                            
                            (tmr_registers(1)(212) and tmr_registers(2)(212)) or                                                       
                            (tmr_registers(0)(212) and tmr_registers(2)(212));                                                         
                                                                                                                                     
        global_tmr_voter(1)(213)  <=    (tmr_registers(0)(213) and tmr_registers(1)(213)) or                                            
                            (tmr_registers(1)(213) and tmr_registers(2)(213)) or                                                       
                            (tmr_registers(0)(213) and tmr_registers(2)(213));                                                         
                                                                                                                                     
        global_tmr_voter(1)(214)  <=    (tmr_registers(0)(214) and tmr_registers(1)(214)) or                                            
                            (tmr_registers(1)(214) and tmr_registers(2)(214)) or                                                       
                            (tmr_registers(0)(214) and tmr_registers(2)(214));                                                         
                                                                                                                                     
        global_tmr_voter(1)(215)  <=    (tmr_registers(0)(215) and tmr_registers(1)(215)) or                                            
                            (tmr_registers(1)(215) and tmr_registers(2)(215)) or                                                       
                            (tmr_registers(0)(215) and tmr_registers(2)(215));                                                         
                                                                                                                                     
        global_tmr_voter(1)(216)  <=    (tmr_registers(0)(216) and tmr_registers(1)(216)) or                                            
                            (tmr_registers(1)(216) and tmr_registers(2)(216)) or                                                       
                            (tmr_registers(0)(216) and tmr_registers(2)(216));                                                         
                                                                                                                                     
        global_tmr_voter(1)(217)  <=    (tmr_registers(0)(217) and tmr_registers(1)(217)) or                                            
                            (tmr_registers(1)(217) and tmr_registers(2)(217)) or                                                       
                            (tmr_registers(0)(217) and tmr_registers(2)(217));                                                         
                                                                                                                                     
        global_tmr_voter(1)(218)  <=    (tmr_registers(0)(218) and tmr_registers(1)(218)) or                                            
                            (tmr_registers(1)(218) and tmr_registers(2)(218)) or                                                       
                            (tmr_registers(0)(218) and tmr_registers(2)(218));                                                         
                                                                                                                                     
        global_tmr_voter(1)(219)  <=    (tmr_registers(0)(219) and tmr_registers(1)(219)) or                                            
                            (tmr_registers(1)(219) and tmr_registers(2)(219)) or                                                       
                            (tmr_registers(0)(219) and tmr_registers(2)(219));                                                         
                                                                                                                                     
        global_tmr_voter(1)(220)  <=    (tmr_registers(0)(220) and tmr_registers(1)(220)) or                                            
                            (tmr_registers(1)(220) and tmr_registers(2)(220)) or                                                       
                            (tmr_registers(0)(220) and tmr_registers(2)(220));                                                         
                                                                                                                                     
        global_tmr_voter(1)(221)  <=    (tmr_registers(0)(221) and tmr_registers(1)(221)) or                                            
                            (tmr_registers(1)(221) and tmr_registers(2)(221)) or                                                       
                            (tmr_registers(0)(221) and tmr_registers(2)(221));                                                         
                                                                                                                                     
        global_tmr_voter(1)(222)  <=    (tmr_registers(0)(222) and tmr_registers(1)(222)) or                                            
                            (tmr_registers(1)(222) and tmr_registers(2)(222)) or                                                       
                            (tmr_registers(0)(222) and tmr_registers(2)(222));                                                         
                                                                                                                                     
        global_tmr_voter(1)(223)  <=    (tmr_registers(0)(223) and tmr_registers(1)(223)) or                                            
                            (tmr_registers(1)(223) and tmr_registers(2)(223)) or                                                       
                            (tmr_registers(0)(223) and tmr_registers(2)(223));                                                         
                                                                                                                                     
        global_tmr_voter(1)(224)  <=    (tmr_registers(0)(224) and tmr_registers(1)(224)) or                                            
                            (tmr_registers(1)(224) and tmr_registers(2)(224)) or                                                       
                            (tmr_registers(0)(224) and tmr_registers(2)(224));                                                         
                                                                                                                                     
        global_tmr_voter(1)(225)  <=    (tmr_registers(0)(225) and tmr_registers(1)(225)) or                                            
                            (tmr_registers(1)(225) and tmr_registers(2)(225)) or                                                       
                            (tmr_registers(0)(225) and tmr_registers(2)(225));                                                         
                                                                                                                                     
        global_tmr_voter(1)(226)  <=    (tmr_registers(0)(226) and tmr_registers(1)(226)) or                                            
                            (tmr_registers(1)(226) and tmr_registers(2)(226)) or                                                       
                            (tmr_registers(0)(226) and tmr_registers(2)(226));                                                         
                                                                                                                                     
        global_tmr_voter(1)(227)  <=    (tmr_registers(0)(227) and tmr_registers(1)(227)) or                                            
                            (tmr_registers(1)(227) and tmr_registers(2)(227)) or                                                       
                            (tmr_registers(0)(227) and tmr_registers(2)(227));                                                         
                                                                                                                                     
        global_tmr_voter(1)(228)  <=    (tmr_registers(0)(228) and tmr_registers(1)(228)) or                                            
                            (tmr_registers(1)(228) and tmr_registers(2)(228)) or                                                       
                            (tmr_registers(0)(228) and tmr_registers(2)(228));                                                         
                                                                                                                                     
        global_tmr_voter(1)(229)  <=    (tmr_registers(0)(229) and tmr_registers(1)(229)) or                                            
                            (tmr_registers(1)(229) and tmr_registers(2)(229)) or                                                       
                            (tmr_registers(0)(229) and tmr_registers(2)(229));                                                         
                                                                                                                                     
        global_tmr_voter(1)(230)  <=    (tmr_registers(0)(230) and tmr_registers(1)(230)) or                                            
                            (tmr_registers(1)(230) and tmr_registers(2)(230)) or                                                       
                            (tmr_registers(0)(230) and tmr_registers(2)(230));                                                         
                                                                                                                                     
        global_tmr_voter(1)(231)  <=    (tmr_registers(0)(231) and tmr_registers(1)(231)) or                                            
                            (tmr_registers(1)(231) and tmr_registers(2)(231)) or                                                       
                            (tmr_registers(0)(231) and tmr_registers(2)(231));                                                         
                                                                                                                                     
        global_tmr_voter(1)(232)  <=    (tmr_registers(0)(232) and tmr_registers(1)(232)) or                                            
                            (tmr_registers(1)(232) and tmr_registers(2)(232)) or                                                       
                            (tmr_registers(0)(232) and tmr_registers(2)(232));                                                         
                                                                                                                                     
        global_tmr_voter(1)(233)  <=    (tmr_registers(0)(233) and tmr_registers(1)(233)) or                                            
                            (tmr_registers(1)(233) and tmr_registers(2)(233)) or                                                       
                            (tmr_registers(0)(233) and tmr_registers(2)(233));                                                         
                                                                                                                                     
        global_tmr_voter(1)(234)  <=    (tmr_registers(0)(234) and tmr_registers(1)(234)) or                                            
                            (tmr_registers(1)(234) and tmr_registers(2)(234)) or                                                       
                            (tmr_registers(0)(234) and tmr_registers(2)(234));                                                         
                                                                                                                                     
        global_tmr_voter(1)(235)  <=    (tmr_registers(0)(235) and tmr_registers(1)(235)) or                                            
                            (tmr_registers(1)(235) and tmr_registers(2)(235)) or                                                       
                            (tmr_registers(0)(235) and tmr_registers(2)(235));                                                         
                                                                                                                                     
        global_tmr_voter(1)(236)  <=    (tmr_registers(0)(236) and tmr_registers(1)(236)) or                                            
                            (tmr_registers(1)(236) and tmr_registers(2)(236)) or                                                       
                            (tmr_registers(0)(236) and tmr_registers(2)(236));                                                         
                                                                                                                                     
        global_tmr_voter(1)(237)  <=    (tmr_registers(0)(237) and tmr_registers(1)(237)) or                                            
                            (tmr_registers(1)(237) and tmr_registers(2)(237)) or                                                       
                            (tmr_registers(0)(237) and tmr_registers(2)(237));                                                         
                                                                                                                                     
        global_tmr_voter(1)(238)  <=    (tmr_registers(0)(238) and tmr_registers(1)(238)) or                                            
                            (tmr_registers(1)(238) and tmr_registers(2)(238)) or                                                       
                            (tmr_registers(0)(238) and tmr_registers(2)(238));                                                         
                                                                                                                                     
        global_tmr_voter(1)(239)  <=    (tmr_registers(0)(239) and tmr_registers(1)(239)) or                                            
                            (tmr_registers(1)(239) and tmr_registers(2)(239)) or                                                       
                            (tmr_registers(0)(239) and tmr_registers(2)(239));                                                         
                                                                                                                                     
        global_tmr_voter(1)(240)  <=    (tmr_registers(0)(240) and tmr_registers(1)(240)) or                                            
                            (tmr_registers(1)(240) and tmr_registers(2)(240)) or                                                       
                            (tmr_registers(0)(240) and tmr_registers(2)(240));                                                         
                                                                                                                                     
        global_tmr_voter(1)(241)  <=    (tmr_registers(0)(241) and tmr_registers(1)(241)) or                                            
                            (tmr_registers(1)(241) and tmr_registers(2)(241)) or                                                       
                            (tmr_registers(0)(241) and tmr_registers(2)(241));                                                         
                                                                                                                                     
        global_tmr_voter(1)(242)  <=    (tmr_registers(0)(242) and tmr_registers(1)(242)) or                                            
                            (tmr_registers(1)(242) and tmr_registers(2)(242)) or                                                       
                            (tmr_registers(0)(242) and tmr_registers(2)(242));                                                         
                                                                                                                                     
        global_tmr_voter(1)(243)  <=    (tmr_registers(0)(243) and tmr_registers(1)(243)) or                                            
                            (tmr_registers(1)(243) and tmr_registers(2)(243)) or                                                       
                            (tmr_registers(0)(243) and tmr_registers(2)(243));                                                         
                                                                                                                                     
        global_tmr_voter(1)(244)  <=    (tmr_registers(0)(244) and tmr_registers(1)(244)) or                                            
                            (tmr_registers(1)(244) and tmr_registers(2)(244)) or                                                       
                            (tmr_registers(0)(244) and tmr_registers(2)(244));                                                         
                                                                                                                                     
        global_tmr_voter(1)(245)  <=    (tmr_registers(0)(245) and tmr_registers(1)(245)) or                                            
                            (tmr_registers(1)(245) and tmr_registers(2)(245)) or                                                       
                            (tmr_registers(0)(245) and tmr_registers(2)(245));                                                         
                                                                                                                                     
        global_tmr_voter(1)(246)  <=    (tmr_registers(0)(246) and tmr_registers(1)(246)) or                                            
                            (tmr_registers(1)(246) and tmr_registers(2)(246)) or                                                       
                            (tmr_registers(0)(246) and tmr_registers(2)(246));                                                         
                                                                                                                                     
        global_tmr_voter(1)(247)  <=    (tmr_registers(0)(247) and tmr_registers(1)(247)) or                                            
                            (tmr_registers(1)(247) and tmr_registers(2)(247)) or                                                       
                            (tmr_registers(0)(247) and tmr_registers(2)(247));                                                         
                                                                                                                                     
        global_tmr_voter(1)(248)  <=    (tmr_registers(0)(248) and tmr_registers(1)(248)) or                                            
                            (tmr_registers(1)(248) and tmr_registers(2)(248)) or                                                       
                            (tmr_registers(0)(248) and tmr_registers(2)(248));                                                         
                                                                                                                                     
        global_tmr_voter(1)(249)  <=    (tmr_registers(0)(249) and tmr_registers(1)(249)) or                                            
                            (tmr_registers(1)(249) and tmr_registers(2)(249)) or                                                       
                            (tmr_registers(0)(249) and tmr_registers(2)(249));                                                         
                                                                                                                                     
        global_tmr_voter(1)(250)  <=    (tmr_registers(0)(250) and tmr_registers(1)(250)) or                                            
                            (tmr_registers(1)(250) and tmr_registers(2)(250)) or                                                       
                            (tmr_registers(0)(250) and tmr_registers(2)(250));                                                         
                                                                                                                                     
        global_tmr_voter(1)(251)  <=    (tmr_registers(0)(251) and tmr_registers(1)(251)) or                                            
                            (tmr_registers(1)(251) and tmr_registers(2)(251)) or                                                       
                            (tmr_registers(0)(251) and tmr_registers(2)(251));                                                         
                                                                                                                                     
        global_tmr_voter(1)(252)  <=    (tmr_registers(0)(252) and tmr_registers(1)(252)) or                                            
                            (tmr_registers(1)(252) and tmr_registers(2)(252)) or                                                       
                            (tmr_registers(0)(252) and tmr_registers(2)(252));                                                         
                                                                                                                                     
        global_tmr_voter(1)(253)  <=    (tmr_registers(0)(253) and tmr_registers(1)(253)) or                                            
                            (tmr_registers(1)(253) and tmr_registers(2)(253)) or                                                       
                            (tmr_registers(0)(253) and tmr_registers(2)(253));                                                         
                                                                                                                                     
        global_tmr_voter(1)(254)  <=    (tmr_registers(0)(254) and tmr_registers(1)(254)) or                                            
                            (tmr_registers(1)(254) and tmr_registers(2)(254)) or                                                       
                            (tmr_registers(0)(254) and tmr_registers(2)(254));                                                         
                                                                                                                                     
        global_tmr_voter(1)(255)  <=    (tmr_registers(0)(255) and tmr_registers(1)(255)) or                                            
                            (tmr_registers(1)(255) and tmr_registers(2)(255)) or                                                       
                            (tmr_registers(0)(255) and tmr_registers(2)(255));                                                         
                                                                                                                                     
        global_tmr_voter(1)(256)  <=    (tmr_registers(0)(256) and tmr_registers(1)(256)) or                                            
                            (tmr_registers(1)(256) and tmr_registers(2)(256)) or                                                       
                            (tmr_registers(0)(256) and tmr_registers(2)(256));                                                         
                                                                                                                                     
        global_tmr_voter(1)(257)  <=    (tmr_registers(0)(257) and tmr_registers(1)(257)) or                                            
                            (tmr_registers(1)(257) and tmr_registers(2)(257)) or                                                       
                            (tmr_registers(0)(257) and tmr_registers(2)(257));                                                         
                                                                                                                                     
        global_tmr_voter(1)(258)  <=    (tmr_registers(0)(258) and tmr_registers(1)(258)) or                                            
                            (tmr_registers(1)(258) and tmr_registers(2)(258)) or                                                       
                            (tmr_registers(0)(258) and tmr_registers(2)(258));                                                         
                                                                                                                                     
        global_tmr_voter(1)(259)  <=    (tmr_registers(0)(259) and tmr_registers(1)(259)) or                                            
                            (tmr_registers(1)(259) and tmr_registers(2)(259)) or                                                       
                            (tmr_registers(0)(259) and tmr_registers(2)(259));                                                         
                                                                                                                                     
        global_tmr_voter(1)(260)  <=    (tmr_registers(0)(260) and tmr_registers(1)(260)) or                                            
                            (tmr_registers(1)(260) and tmr_registers(2)(260)) or                                                       
                            (tmr_registers(0)(260) and tmr_registers(2)(260));                                                         
                                                                                                                                     
        global_tmr_voter(1)(261)  <=    (tmr_registers(0)(261) and tmr_registers(1)(261)) or                                            
                            (tmr_registers(1)(261) and tmr_registers(2)(261)) or                                                       
                            (tmr_registers(0)(261) and tmr_registers(2)(261));                                                         
                                                                                                                                     
        global_tmr_voter(1)(262)  <=    (tmr_registers(0)(262) and tmr_registers(1)(262)) or                                            
                            (tmr_registers(1)(262) and tmr_registers(2)(262)) or                                                       
                            (tmr_registers(0)(262) and tmr_registers(2)(262));                                                         
                                                                                                                                     
        global_tmr_voter(1)(263)  <=    (tmr_registers(0)(263) and tmr_registers(1)(263)) or                                            
                            (tmr_registers(1)(263) and tmr_registers(2)(263)) or                                                       
                            (tmr_registers(0)(263) and tmr_registers(2)(263));                                                         
                                                                                                                                     
        global_tmr_voter(1)(264)  <=    (tmr_registers(0)(264) and tmr_registers(1)(264)) or                                            
                            (tmr_registers(1)(264) and tmr_registers(2)(264)) or                                                       
                            (tmr_registers(0)(264) and tmr_registers(2)(264));                                                         
                                                                                                                                     
        global_tmr_voter(1)(265)  <=    (tmr_registers(0)(265) and tmr_registers(1)(265)) or                                            
                            (tmr_registers(1)(265) and tmr_registers(2)(265)) or                                                       
                            (tmr_registers(0)(265) and tmr_registers(2)(265));                                                         
                                                                                                                                     
        global_tmr_voter(1)(266)  <=    (tmr_registers(0)(266) and tmr_registers(1)(266)) or                                            
                            (tmr_registers(1)(266) and tmr_registers(2)(266)) or                                                       
                            (tmr_registers(0)(266) and tmr_registers(2)(266));                                                         
                                                                                                                                     
        global_tmr_voter(1)(267)  <=    (tmr_registers(0)(267) and tmr_registers(1)(267)) or                                            
                            (tmr_registers(1)(267) and tmr_registers(2)(267)) or                                                       
                            (tmr_registers(0)(267) and tmr_registers(2)(267));                                                         
                                                                                                                                     
        global_tmr_voter(1)(268)  <=    (tmr_registers(0)(268) and tmr_registers(1)(268)) or                                            
                            (tmr_registers(1)(268) and tmr_registers(2)(268)) or                                                       
                            (tmr_registers(0)(268) and tmr_registers(2)(268));                                                         
                                                                                                                                     
        global_tmr_voter(1)(269)  <=    (tmr_registers(0)(269) and tmr_registers(1)(269)) or                                            
                            (tmr_registers(1)(269) and tmr_registers(2)(269)) or                                                       
                            (tmr_registers(0)(269) and tmr_registers(2)(269));                                                         
                                                                                                                                     
        global_tmr_voter(1)(270)  <=    (tmr_registers(0)(270) and tmr_registers(1)(270)) or                                            
                            (tmr_registers(1)(270) and tmr_registers(2)(270)) or                                                       
                            (tmr_registers(0)(270) and tmr_registers(2)(270));                                                         
                                                                                                                                     
        global_tmr_voter(1)(271)  <=    (tmr_registers(0)(271) and tmr_registers(1)(271)) or                                            
                            (tmr_registers(1)(271) and tmr_registers(2)(271)) or                                                       
                            (tmr_registers(0)(271) and tmr_registers(2)(271));                                                         
                                                                                                                                     
        global_tmr_voter(1)(272)  <=    (tmr_registers(0)(272) and tmr_registers(1)(272)) or                                            
                            (tmr_registers(1)(272) and tmr_registers(2)(272)) or                                                       
                            (tmr_registers(0)(272) and tmr_registers(2)(272));                                                         
                                                                                                                                     
        global_tmr_voter(1)(273)  <=    (tmr_registers(0)(273) and tmr_registers(1)(273)) or                                            
                            (tmr_registers(1)(273) and tmr_registers(2)(273)) or                                                       
                            (tmr_registers(0)(273) and tmr_registers(2)(273));                                                         
                                                                                                                                     
        global_tmr_voter(1)(274)  <=    (tmr_registers(0)(274) and tmr_registers(1)(274)) or                                            
                            (tmr_registers(1)(274) and tmr_registers(2)(274)) or                                                       
                            (tmr_registers(0)(274) and tmr_registers(2)(274));                                                         
                                                                                                                                     
        global_tmr_voter(1)(275)  <=    (tmr_registers(0)(275) and tmr_registers(1)(275)) or                                            
                            (tmr_registers(1)(275) and tmr_registers(2)(275)) or                                                       
                            (tmr_registers(0)(275) and tmr_registers(2)(275));                                                         
                                                                                                                                     
        global_tmr_voter(1)(276)  <=    (tmr_registers(0)(276) and tmr_registers(1)(276)) or                                            
                            (tmr_registers(1)(276) and tmr_registers(2)(276)) or                                                       
                            (tmr_registers(0)(276) and tmr_registers(2)(276));                                                         
                                                                                                                                     
        global_tmr_voter(1)(277)  <=    (tmr_registers(0)(277) and tmr_registers(1)(277)) or                                            
                            (tmr_registers(1)(277) and tmr_registers(2)(277)) or                                                       
                            (tmr_registers(0)(277) and tmr_registers(2)(277));                                                         
                                                                                                                                     
        global_tmr_voter(1)(278)  <=    (tmr_registers(0)(278) and tmr_registers(1)(278)) or                                            
                            (tmr_registers(1)(278) and tmr_registers(2)(278)) or                                                       
                            (tmr_registers(0)(278) and tmr_registers(2)(278));                                                         
                                                                                                                                     
        global_tmr_voter(1)(279)  <=    (tmr_registers(0)(279) and tmr_registers(1)(279)) or                                            
                            (tmr_registers(1)(279) and tmr_registers(2)(279)) or                                                       
                            (tmr_registers(0)(279) and tmr_registers(2)(279));                                                         
                                                                                                                                     
        global_tmr_voter(1)(280)  <=    (tmr_registers(0)(280) and tmr_registers(1)(280)) or                                            
                            (tmr_registers(1)(280) and tmr_registers(2)(280)) or                                                       
                            (tmr_registers(0)(280) and tmr_registers(2)(280));                                                         
                                                                                                                                     
        global_tmr_voter(1)(281)  <=    (tmr_registers(0)(281) and tmr_registers(1)(281)) or                                            
                            (tmr_registers(1)(281) and tmr_registers(2)(281)) or                                                       
                            (tmr_registers(0)(281) and tmr_registers(2)(281));                                                         
                                                                                                                                     
        global_tmr_voter(1)(282)  <=    (tmr_registers(0)(282) and tmr_registers(1)(282)) or                                            
                            (tmr_registers(1)(282) and tmr_registers(2)(282)) or                                                       
                            (tmr_registers(0)(282) and tmr_registers(2)(282));                                                         
                                                                                                                                     
        global_tmr_voter(1)(283)  <=    (tmr_registers(0)(283) and tmr_registers(1)(283)) or                                            
                            (tmr_registers(1)(283) and tmr_registers(2)(283)) or                                                       
                            (tmr_registers(0)(283) and tmr_registers(2)(283));                                                         
                                                                                                                                     
        global_tmr_voter(1)(284)  <=    (tmr_registers(0)(284) and tmr_registers(1)(284)) or                                            
                            (tmr_registers(1)(284) and tmr_registers(2)(284)) or                                                       
                            (tmr_registers(0)(284) and tmr_registers(2)(284));                                                         
                                                                                                                                     
        global_tmr_voter(1)(285)  <=    (tmr_registers(0)(285) and tmr_registers(1)(285)) or                                            
                            (tmr_registers(1)(285) and tmr_registers(2)(285)) or                                                       
                            (tmr_registers(0)(285) and tmr_registers(2)(285));                                                         
                                                                                                                                     
        global_tmr_voter(1)(286)  <=    (tmr_registers(0)(286) and tmr_registers(1)(286)) or                                            
                            (tmr_registers(1)(286) and tmr_registers(2)(286)) or                                                       
                            (tmr_registers(0)(286) and tmr_registers(2)(286));                                                         
                                                                                                                                     
        global_tmr_voter(1)(287)  <=    (tmr_registers(0)(287) and tmr_registers(1)(287)) or                                            
                            (tmr_registers(1)(287) and tmr_registers(2)(287)) or                                                       
                            (tmr_registers(0)(287) and tmr_registers(2)(287));                                                         
                                                                                                                                     
        global_tmr_voter(1)(288)  <=    (tmr_registers(0)(288) and tmr_registers(1)(288)) or                                            
                            (tmr_registers(1)(288) and tmr_registers(2)(288)) or                                                       
                            (tmr_registers(0)(288) and tmr_registers(2)(288));                                                         
                                                                                                                                     
        global_tmr_voter(1)(289)  <=    (tmr_registers(0)(289) and tmr_registers(1)(289)) or                                            
                            (tmr_registers(1)(289) and tmr_registers(2)(289)) or                                                       
                            (tmr_registers(0)(289) and tmr_registers(2)(289));                                                         
                                                                                                                                     
        global_tmr_voter(1)(290)  <=    (tmr_registers(0)(290) and tmr_registers(1)(290)) or                                            
                            (tmr_registers(1)(290) and tmr_registers(2)(290)) or                                                       
                            (tmr_registers(0)(290) and tmr_registers(2)(290));                                                         
                                                                                                                                     
        global_tmr_voter(1)(291)  <=    (tmr_registers(0)(291) and tmr_registers(1)(291)) or                                            
                            (tmr_registers(1)(291) and tmr_registers(2)(291)) or                                                       
                            (tmr_registers(0)(291) and tmr_registers(2)(291));                                                         
                                                                                                                                     
        global_tmr_voter(1)(292)  <=    (tmr_registers(0)(292) and tmr_registers(1)(292)) or                                            
                            (tmr_registers(1)(292) and tmr_registers(2)(292)) or                                                       
                            (tmr_registers(0)(292) and tmr_registers(2)(292));                                                         
                                                                                                                                     
        global_tmr_voter(1)(293)  <=    (tmr_registers(0)(293) and tmr_registers(1)(293)) or                                            
                            (tmr_registers(1)(293) and tmr_registers(2)(293)) or                                                       
                            (tmr_registers(0)(293) and tmr_registers(2)(293));                                                         
                                                                                                                                     
        global_tmr_voter(1)(294)  <=    (tmr_registers(0)(294) and tmr_registers(1)(294)) or                                            
                            (tmr_registers(1)(294) and tmr_registers(2)(294)) or                                                       
                            (tmr_registers(0)(294) and tmr_registers(2)(294));                                                         
                                                                                                                                     
        global_tmr_voter(1)(295)  <=    (tmr_registers(0)(295) and tmr_registers(1)(295)) or                                            
                            (tmr_registers(1)(295) and tmr_registers(2)(295)) or                                                       
                            (tmr_registers(0)(295) and tmr_registers(2)(295));                                                         
                                                                                                                                     
        global_tmr_voter(1)(296)  <=    (tmr_registers(0)(296) and tmr_registers(1)(296)) or                                            
                            (tmr_registers(1)(296) and tmr_registers(2)(296)) or                                                       
                            (tmr_registers(0)(296) and tmr_registers(2)(296));                                                         
                                                                                                                                     
        global_tmr_voter(1)(297)  <=    (tmr_registers(0)(297) and tmr_registers(1)(297)) or                                            
                            (tmr_registers(1)(297) and tmr_registers(2)(297)) or                                                       
                            (tmr_registers(0)(297) and tmr_registers(2)(297));                                                         
                                                                                                                                     
        global_tmr_voter(1)(298)  <=    (tmr_registers(0)(298) and tmr_registers(1)(298)) or                                            
                            (tmr_registers(1)(298) and tmr_registers(2)(298)) or                                                       
                            (tmr_registers(0)(298) and tmr_registers(2)(298));                                                         
                                                                                                                                     
        global_tmr_voter(1)(299)  <=    (tmr_registers(0)(299) and tmr_registers(1)(299)) or                                            
                            (tmr_registers(1)(299) and tmr_registers(2)(299)) or                                                       
                            (tmr_registers(0)(299) and tmr_registers(2)(299));                                                         
                                                                                                                                     
        global_tmr_voter(1)(300)  <=    (tmr_registers(0)(300) and tmr_registers(1)(300)) or                                            
                            (tmr_registers(1)(300) and tmr_registers(2)(300)) or                                                       
                            (tmr_registers(0)(300) and tmr_registers(2)(300));                                                         
                                                                                                                                     
        global_tmr_voter(1)(301)  <=    (tmr_registers(0)(301) and tmr_registers(1)(301)) or                                            
                            (tmr_registers(1)(301) and tmr_registers(2)(301)) or                                                       
                            (tmr_registers(0)(301) and tmr_registers(2)(301));                                                         
                                                                                                                                     
        global_tmr_voter(1)(302)  <=    (tmr_registers(0)(302) and tmr_registers(1)(302)) or                                            
                            (tmr_registers(1)(302) and tmr_registers(2)(302)) or                                                       
                            (tmr_registers(0)(302) and tmr_registers(2)(302));                                                         
                                                                                                                                     
        global_tmr_voter(1)(303)  <=    (tmr_registers(0)(303) and tmr_registers(1)(303)) or                                            
                            (tmr_registers(1)(303) and tmr_registers(2)(303)) or                                                       
                            (tmr_registers(0)(303) and tmr_registers(2)(303));                                                         
                                                                                                                                     
        global_tmr_voter(1)(304)  <=    (tmr_registers(0)(304) and tmr_registers(1)(304)) or                                            
                            (tmr_registers(1)(304) and tmr_registers(2)(304)) or                                                       
                            (tmr_registers(0)(304) and tmr_registers(2)(304));                                                         
                                                                                                                                     
        global_tmr_voter(1)(305)  <=    (tmr_registers(0)(305) and tmr_registers(1)(305)) or                                            
                            (tmr_registers(1)(305) and tmr_registers(2)(305)) or                                                       
                            (tmr_registers(0)(305) and tmr_registers(2)(305));                                                         
                                                                                                                                     
        global_tmr_voter(1)(306)  <=    (tmr_registers(0)(306) and tmr_registers(1)(306)) or                                            
                            (tmr_registers(1)(306) and tmr_registers(2)(306)) or                                                       
                            (tmr_registers(0)(306) and tmr_registers(2)(306));                                                         
                                                                                                                                     
        global_tmr_voter(1)(307)  <=    (tmr_registers(0)(307) and tmr_registers(1)(307)) or                                            
                            (tmr_registers(1)(307) and tmr_registers(2)(307)) or                                                       
                            (tmr_registers(0)(307) and tmr_registers(2)(307));                                                         
                                                                                                                                     
        global_tmr_voter(1)(308)  <=    (tmr_registers(0)(308) and tmr_registers(1)(308)) or                                            
                            (tmr_registers(1)(308) and tmr_registers(2)(308)) or                                                       
                            (tmr_registers(0)(308) and tmr_registers(2)(308));                                                         
                                                                                                                                     
        global_tmr_voter(1)(309)  <=    (tmr_registers(0)(309) and tmr_registers(1)(309)) or                                            
                            (tmr_registers(1)(309) and tmr_registers(2)(309)) or                                                       
                            (tmr_registers(0)(309) and tmr_registers(2)(309));                                                         
                                                                                                                                     
        global_tmr_voter(1)(310)  <=    (tmr_registers(0)(310) and tmr_registers(1)(310)) or                                            
                            (tmr_registers(1)(310) and tmr_registers(2)(310)) or                                                       
                            (tmr_registers(0)(310) and tmr_registers(2)(310));                                                         
                                                                                                                                     
        global_tmr_voter(1)(311)  <=    (tmr_registers(0)(311) and tmr_registers(1)(311)) or                                            
                            (tmr_registers(1)(311) and tmr_registers(2)(311)) or                                                       
                            (tmr_registers(0)(311) and tmr_registers(2)(311));                                                         
                                                                                                                                     
        global_tmr_voter(1)(312)  <=    (tmr_registers(0)(312) and tmr_registers(1)(312)) or                                            
                            (tmr_registers(1)(312) and tmr_registers(2)(312)) or                                                       
                            (tmr_registers(0)(312) and tmr_registers(2)(312));                                                         
                                                                                                                                     
        global_tmr_voter(1)(313)  <=    (tmr_registers(0)(313) and tmr_registers(1)(313)) or                                            
                            (tmr_registers(1)(313) and tmr_registers(2)(313)) or                                                       
                            (tmr_registers(0)(313) and tmr_registers(2)(313));                                                         
                                                                                                                                     
        global_tmr_voter(1)(314)  <=    (tmr_registers(0)(314) and tmr_registers(1)(314)) or                                            
                            (tmr_registers(1)(314) and tmr_registers(2)(314)) or                                                       
                            (tmr_registers(0)(314) and tmr_registers(2)(314));                                                         
                                                                                                                                     
        global_tmr_voter(1)(315)  <=    (tmr_registers(0)(315) and tmr_registers(1)(315)) or                                            
                            (tmr_registers(1)(315) and tmr_registers(2)(315)) or                                                       
                            (tmr_registers(0)(315) and tmr_registers(2)(315));                                                         
                                                                                                                                     
        global_tmr_voter(1)(316)  <=    (tmr_registers(0)(316) and tmr_registers(1)(316)) or                                            
                            (tmr_registers(1)(316) and tmr_registers(2)(316)) or                                                       
                            (tmr_registers(0)(316) and tmr_registers(2)(316));                                                         
                                                                                                                                     
        global_tmr_voter(1)(317)  <=    (tmr_registers(0)(317) and tmr_registers(1)(317)) or                                            
                            (tmr_registers(1)(317) and tmr_registers(2)(317)) or                                                       
                            (tmr_registers(0)(317) and tmr_registers(2)(317));                                                         
                                                                                                                                     
        global_tmr_voter(1)(318)  <=    (tmr_registers(0)(318) and tmr_registers(1)(318)) or                                            
                            (tmr_registers(1)(318) and tmr_registers(2)(318)) or                                                       
                            (tmr_registers(0)(318) and tmr_registers(2)(318));                                                         
                                                                                                                                     
        global_tmr_voter(1)(319)  <=    (tmr_registers(0)(319) and tmr_registers(1)(319)) or                                            
                            (tmr_registers(1)(319) and tmr_registers(2)(319)) or                                                       
                            (tmr_registers(0)(319) and tmr_registers(2)(319));                                                         
                                                                                                                                     
        global_tmr_voter(1)(320)  <=    (tmr_registers(0)(320) and tmr_registers(1)(320)) or                                            
                            (tmr_registers(1)(320) and tmr_registers(2)(320)) or                                                       
                            (tmr_registers(0)(320) and tmr_registers(2)(320));                                                         
                                                                                                                                     
        global_tmr_voter(1)(321)  <=    (tmr_registers(0)(321) and tmr_registers(1)(321)) or                                            
                            (tmr_registers(1)(321) and tmr_registers(2)(321)) or                                                       
                            (tmr_registers(0)(321) and tmr_registers(2)(321));                                                         
                                                                                                                                     
        global_tmr_voter(1)(322)  <=    (tmr_registers(0)(322) and tmr_registers(1)(322)) or                                            
                            (tmr_registers(1)(322) and tmr_registers(2)(322)) or                                                       
                            (tmr_registers(0)(322) and tmr_registers(2)(322));                                                         
                                                                                                                                     
        global_tmr_voter(1)(323)  <=    (tmr_registers(0)(323) and tmr_registers(1)(323)) or                                            
                            (tmr_registers(1)(323) and tmr_registers(2)(323)) or                                                       
                            (tmr_registers(0)(323) and tmr_registers(2)(323));                                                         
                                                                                                                                     
        global_tmr_voter(1)(324)  <=    (tmr_registers(0)(324) and tmr_registers(1)(324)) or                                            
                            (tmr_registers(1)(324) and tmr_registers(2)(324)) or                                                       
                            (tmr_registers(0)(324) and tmr_registers(2)(324));                                                         
                                                                                                                                     
        global_tmr_voter(1)(325)  <=    (tmr_registers(0)(325) and tmr_registers(1)(325)) or                                            
                            (tmr_registers(1)(325) and tmr_registers(2)(325)) or                                                       
                            (tmr_registers(0)(325) and tmr_registers(2)(325));                                                         
                                                                                                                                     
        global_tmr_voter(1)(326)  <=    (tmr_registers(0)(326) and tmr_registers(1)(326)) or                                            
                            (tmr_registers(1)(326) and tmr_registers(2)(326)) or                                                       
                            (tmr_registers(0)(326) and tmr_registers(2)(326));                                                         
                                                                                                                                     
        global_tmr_voter(1)(327)  <=    (tmr_registers(0)(327) and tmr_registers(1)(327)) or                                            
                            (tmr_registers(1)(327) and tmr_registers(2)(327)) or                                                       
                            (tmr_registers(0)(327) and tmr_registers(2)(327));                                                         
                                                                                                                                     
        global_tmr_voter(1)(328)  <=    (tmr_registers(0)(328) and tmr_registers(1)(328)) or                                            
                            (tmr_registers(1)(328) and tmr_registers(2)(328)) or                                                       
                            (tmr_registers(0)(328) and tmr_registers(2)(328));                                                         
                                                                                                                                     
        global_tmr_voter(1)(329)  <=    (tmr_registers(0)(329) and tmr_registers(1)(329)) or                                            
                            (tmr_registers(1)(329) and tmr_registers(2)(329)) or                                                       
                            (tmr_registers(0)(329) and tmr_registers(2)(329));                                                         
                                                                                                                                     
        global_tmr_voter(1)(330)  <=    (tmr_registers(0)(330) and tmr_registers(1)(330)) or                                            
                            (tmr_registers(1)(330) and tmr_registers(2)(330)) or                                                       
                            (tmr_registers(0)(330) and tmr_registers(2)(330));                                                         
                                                                                                                                     
        global_tmr_voter(1)(331)  <=    (tmr_registers(0)(331) and tmr_registers(1)(331)) or                                            
                            (tmr_registers(1)(331) and tmr_registers(2)(331)) or                                                       
                            (tmr_registers(0)(331) and tmr_registers(2)(331));                                                         
                                                                                                                                     
        global_tmr_voter(1)(332)  <=    (tmr_registers(0)(332) and tmr_registers(1)(332)) or                                            
                            (tmr_registers(1)(332) and tmr_registers(2)(332)) or                                                       
                            (tmr_registers(0)(332) and tmr_registers(2)(332));                                                         
                                                                                                                                     
        global_tmr_voter(1)(333)  <=    (tmr_registers(0)(333) and tmr_registers(1)(333)) or                                            
                            (tmr_registers(1)(333) and tmr_registers(2)(333)) or                                                       
                            (tmr_registers(0)(333) and tmr_registers(2)(333));                                                         
                                                                                                                                     
        global_tmr_voter(1)(334)  <=    (tmr_registers(0)(334) and tmr_registers(1)(334)) or                                            
                            (tmr_registers(1)(334) and tmr_registers(2)(334)) or                                                       
                            (tmr_registers(0)(334) and tmr_registers(2)(334));                                                         
                                                                                                                                     
        global_tmr_voter(1)(335)  <=    (tmr_registers(0)(335) and tmr_registers(1)(335)) or                                            
                            (tmr_registers(1)(335) and tmr_registers(2)(335)) or                                                       
                            (tmr_registers(0)(335) and tmr_registers(2)(335));                                                         
                                                                                                                                     
        global_tmr_voter(1)(336)  <=    (tmr_registers(0)(336) and tmr_registers(1)(336)) or                                            
                            (tmr_registers(1)(336) and tmr_registers(2)(336)) or                                                       
                            (tmr_registers(0)(336) and tmr_registers(2)(336));                                                         
                                                                                                                                     
        global_tmr_voter(1)(337)  <=    (tmr_registers(0)(337) and tmr_registers(1)(337)) or                                            
                            (tmr_registers(1)(337) and tmr_registers(2)(337)) or                                                       
                            (tmr_registers(0)(337) and tmr_registers(2)(337));                                                         
                                                                                                                                     
        global_tmr_voter(1)(338)  <=    (tmr_registers(0)(338) and tmr_registers(1)(338)) or                                            
                            (tmr_registers(1)(338) and tmr_registers(2)(338)) or                                                       
                            (tmr_registers(0)(338) and tmr_registers(2)(338));                                                         
                                                                                                                                     
        global_tmr_voter(1)(339)  <=    (tmr_registers(0)(339) and tmr_registers(1)(339)) or                                            
                            (tmr_registers(1)(339) and tmr_registers(2)(339)) or                                                       
                            (tmr_registers(0)(339) and tmr_registers(2)(339));                                                         
                                                                                                                                     
        global_tmr_voter(1)(340)  <=    (tmr_registers(0)(340) and tmr_registers(1)(340)) or                                            
                            (tmr_registers(1)(340) and tmr_registers(2)(340)) or                                                       
                            (tmr_registers(0)(340) and tmr_registers(2)(340));                                                         
                                                                                                                                     
        global_tmr_voter(1)(341)  <=    (tmr_registers(0)(341) and tmr_registers(1)(341)) or                                            
                            (tmr_registers(1)(341) and tmr_registers(2)(341)) or                                                       
                            (tmr_registers(0)(341) and tmr_registers(2)(341));                                                         
                                                                                                                                     
        global_tmr_voter(1)(342)  <=    (tmr_registers(0)(342) and tmr_registers(1)(342)) or                                            
                            (tmr_registers(1)(342) and tmr_registers(2)(342)) or                                                       
                            (tmr_registers(0)(342) and tmr_registers(2)(342));                                                         
                                                                                                                                     
        global_tmr_voter(1)(343)  <=    (tmr_registers(0)(343) and tmr_registers(1)(343)) or                                            
                            (tmr_registers(1)(343) and tmr_registers(2)(343)) or                                                       
                            (tmr_registers(0)(343) and tmr_registers(2)(343));                                                         
                                                                                                                                     
        global_tmr_voter(1)(344)  <=    (tmr_registers(0)(344) and tmr_registers(1)(344)) or                                            
                            (tmr_registers(1)(344) and tmr_registers(2)(344)) or                                                       
                            (tmr_registers(0)(344) and tmr_registers(2)(344));                                                         
                                                                                                                                     
        global_tmr_voter(1)(345)  <=    (tmr_registers(0)(345) and tmr_registers(1)(345)) or                                            
                            (tmr_registers(1)(345) and tmr_registers(2)(345)) or                                                       
                            (tmr_registers(0)(345) and tmr_registers(2)(345));                                                         
                                                                                                                                     
        global_tmr_voter(1)(346)  <=    (tmr_registers(0)(346) and tmr_registers(1)(346)) or                                            
                            (tmr_registers(1)(346) and tmr_registers(2)(346)) or                                                       
                            (tmr_registers(0)(346) and tmr_registers(2)(346));                                                         
                                                                                                                                     
        global_tmr_voter(1)(347)  <=    (tmr_registers(0)(347) and tmr_registers(1)(347)) or                                            
                            (tmr_registers(1)(347) and tmr_registers(2)(347)) or                                                       
                            (tmr_registers(0)(347) and tmr_registers(2)(347));                                                         
                                                                                                                                     
        global_tmr_voter(1)(348)  <=    (tmr_registers(0)(348) and tmr_registers(1)(348)) or                                            
                            (tmr_registers(1)(348) and tmr_registers(2)(348)) or                                                       
                            (tmr_registers(0)(348) and tmr_registers(2)(348));                                                         
                                                                                                                                     
        global_tmr_voter(1)(349)  <=    (tmr_registers(0)(349) and tmr_registers(1)(349)) or                                            
                            (tmr_registers(1)(349) and tmr_registers(2)(349)) or                                                       
                            (tmr_registers(0)(349) and tmr_registers(2)(349));                                                         
                                                                                                                                     
        global_tmr_voter(1)(350)  <=    (tmr_registers(0)(350) and tmr_registers(1)(350)) or                                            
                            (tmr_registers(1)(350) and tmr_registers(2)(350)) or                                                       
                            (tmr_registers(0)(350) and tmr_registers(2)(350));                                                         
                                                                                                                                     
        global_tmr_voter(1)(351)  <=    (tmr_registers(0)(351) and tmr_registers(1)(351)) or                                            
                            (tmr_registers(1)(351) and tmr_registers(2)(351)) or                                                       
                            (tmr_registers(0)(351) and tmr_registers(2)(351));                                                         
                                                                                                                                     
        global_tmr_voter(1)(352)  <=    (tmr_registers(0)(352) and tmr_registers(1)(352)) or                                            
                            (tmr_registers(1)(352) and tmr_registers(2)(352)) or                                                       
                            (tmr_registers(0)(352) and tmr_registers(2)(352));                                                         
                                                                                                                                     
        global_tmr_voter(1)(353)  <=    (tmr_registers(0)(353) and tmr_registers(1)(353)) or                                            
                            (tmr_registers(1)(353) and tmr_registers(2)(353)) or                                                       
                            (tmr_registers(0)(353) and tmr_registers(2)(353));                                                         
                                                                                                                                     
        global_tmr_voter(1)(354)  <=    (tmr_registers(0)(354) and tmr_registers(1)(354)) or                                            
                            (tmr_registers(1)(354) and tmr_registers(2)(354)) or                                                       
                            (tmr_registers(0)(354) and tmr_registers(2)(354));                                                         
                                                                                                                                     
        global_tmr_voter(1)(355)  <=    (tmr_registers(0)(355) and tmr_registers(1)(355)) or                                            
                            (tmr_registers(1)(355) and tmr_registers(2)(355)) or                                                       
                            (tmr_registers(0)(355) and tmr_registers(2)(355));                                                         
                                                                                                                                     
        global_tmr_voter(1)(356)  <=    (tmr_registers(0)(356) and tmr_registers(1)(356)) or                                            
                            (tmr_registers(1)(356) and tmr_registers(2)(356)) or                                                       
                            (tmr_registers(0)(356) and tmr_registers(2)(356));                                                         
                                                                                                                                     
        global_tmr_voter(1)(357)  <=    (tmr_registers(0)(357) and tmr_registers(1)(357)) or                                            
                            (tmr_registers(1)(357) and tmr_registers(2)(357)) or                                                       
                            (tmr_registers(0)(357) and tmr_registers(2)(357));                                                         
                                                                                                                                     
        global_tmr_voter(1)(358)  <=    (tmr_registers(0)(358) and tmr_registers(1)(358)) or                                            
                            (tmr_registers(1)(358) and tmr_registers(2)(358)) or                                                       
                            (tmr_registers(0)(358) and tmr_registers(2)(358));                                                         
                                                                                                                                     
        global_tmr_voter(1)(359)  <=    (tmr_registers(0)(359) and tmr_registers(1)(359)) or                                            
                            (tmr_registers(1)(359) and tmr_registers(2)(359)) or                                                       
                            (tmr_registers(0)(359) and tmr_registers(2)(359));                                                         
                                                                                                                                     
        global_tmr_voter(1)(360)  <=    (tmr_registers(0)(360) and tmr_registers(1)(360)) or                                            
                            (tmr_registers(1)(360) and tmr_registers(2)(360)) or                                                       
                            (tmr_registers(0)(360) and tmr_registers(2)(360));                                                         
                                                                                                                                     
        global_tmr_voter(1)(361)  <=    (tmr_registers(0)(361) and tmr_registers(1)(361)) or                                            
                            (tmr_registers(1)(361) and tmr_registers(2)(361)) or                                                       
                            (tmr_registers(0)(361) and tmr_registers(2)(361));                                                         
                                                                                                                                     
        global_tmr_voter(1)(362)  <=    (tmr_registers(0)(362) and tmr_registers(1)(362)) or                                            
                            (tmr_registers(1)(362) and tmr_registers(2)(362)) or                                                       
                            (tmr_registers(0)(362) and tmr_registers(2)(362));                                                         
                                                                                                                                     
        global_tmr_voter(1)(363)  <=    (tmr_registers(0)(363) and tmr_registers(1)(363)) or                                            
                            (tmr_registers(1)(363) and tmr_registers(2)(363)) or                                                       
                            (tmr_registers(0)(363) and tmr_registers(2)(363));                                                         
                                                                                                                                     
        global_tmr_voter(1)(364)  <=    (tmr_registers(0)(364) and tmr_registers(1)(364)) or                                            
                            (tmr_registers(1)(364) and tmr_registers(2)(364)) or                                                       
                            (tmr_registers(0)(364) and tmr_registers(2)(364));                                                         
                                                                                                                                     
        global_tmr_voter(1)(365)  <=    (tmr_registers(0)(365) and tmr_registers(1)(365)) or                                            
                            (tmr_registers(1)(365) and tmr_registers(2)(365)) or                                                       
                            (tmr_registers(0)(365) and tmr_registers(2)(365));                                                         
                                                                                                                                     
        global_tmr_voter(1)(366)  <=    (tmr_registers(0)(366) and tmr_registers(1)(366)) or                                            
                            (tmr_registers(1)(366) and tmr_registers(2)(366)) or                                                       
                            (tmr_registers(0)(366) and tmr_registers(2)(366));                                                         
                                                                                                                                     
        global_tmr_voter(1)(367)  <=    (tmr_registers(0)(367) and tmr_registers(1)(367)) or                                            
                            (tmr_registers(1)(367) and tmr_registers(2)(367)) or                                                       
                            (tmr_registers(0)(367) and tmr_registers(2)(367));                                                         
                                                                                                                                     
        global_tmr_voter(1)(368)  <=    (tmr_registers(0)(368) and tmr_registers(1)(368)) or                                            
                            (tmr_registers(1)(368) and tmr_registers(2)(368)) or                                                       
                            (tmr_registers(0)(368) and tmr_registers(2)(368));                                                         
                                                                                                                                     
        global_tmr_voter(1)(369)  <=    (tmr_registers(0)(369) and tmr_registers(1)(369)) or                                            
                            (tmr_registers(1)(369) and tmr_registers(2)(369)) or                                                       
                            (tmr_registers(0)(369) and tmr_registers(2)(369));                                                         
                                                                                                                                     
        global_tmr_voter(1)(370)  <=    (tmr_registers(0)(370) and tmr_registers(1)(370)) or                                            
                            (tmr_registers(1)(370) and tmr_registers(2)(370)) or                                                       
                            (tmr_registers(0)(370) and tmr_registers(2)(370));                                                         
                                                                                                                                     
        global_tmr_voter(1)(371)  <=    (tmr_registers(0)(371) and tmr_registers(1)(371)) or                                            
                            (tmr_registers(1)(371) and tmr_registers(2)(371)) or                                                       
                            (tmr_registers(0)(371) and tmr_registers(2)(371));                                                         
                                                                                                                                     
        global_tmr_voter(1)(372)  <=    (tmr_registers(0)(372) and tmr_registers(1)(372)) or                                            
                            (tmr_registers(1)(372) and tmr_registers(2)(372)) or                                                       
                            (tmr_registers(0)(372) and tmr_registers(2)(372));                                                         
                                                                                                                                     
        global_tmr_voter(1)(373)  <=    (tmr_registers(0)(373) and tmr_registers(1)(373)) or                                            
                            (tmr_registers(1)(373) and tmr_registers(2)(373)) or                                                       
                            (tmr_registers(0)(373) and tmr_registers(2)(373));                                                         
                                                                                                                                     
        global_tmr_voter(1)(374)  <=    (tmr_registers(0)(374) and tmr_registers(1)(374)) or                                            
                            (tmr_registers(1)(374) and tmr_registers(2)(374)) or                                                       
                            (tmr_registers(0)(374) and tmr_registers(2)(374));                                                         
                                                                                                                                     
        global_tmr_voter(1)(375)  <=    (tmr_registers(0)(375) and tmr_registers(1)(375)) or                                            
                            (tmr_registers(1)(375) and tmr_registers(2)(375)) or                                                       
                            (tmr_registers(0)(375) and tmr_registers(2)(375));                                                         
                                                                                                                                     
        global_tmr_voter(1)(376)  <=    (tmr_registers(0)(376) and tmr_registers(1)(376)) or                                            
                            (tmr_registers(1)(376) and tmr_registers(2)(376)) or                                                       
                            (tmr_registers(0)(376) and tmr_registers(2)(376));                                                         
                                                                                                                                     
        global_tmr_voter(1)(377)  <=    (tmr_registers(0)(377) and tmr_registers(1)(377)) or                                            
                            (tmr_registers(1)(377) and tmr_registers(2)(377)) or                                                       
                            (tmr_registers(0)(377) and tmr_registers(2)(377));                                                         
                                                                                                                                     
        global_tmr_voter(1)(378)  <=    (tmr_registers(0)(378) and tmr_registers(1)(378)) or                                            
                            (tmr_registers(1)(378) and tmr_registers(2)(378)) or                                                       
                            (tmr_registers(0)(378) and tmr_registers(2)(378));                                                         
                                                                                                                                     
        global_tmr_voter(1)(379)  <=    (tmr_registers(0)(379) and tmr_registers(1)(379)) or                                            
                            (tmr_registers(1)(379) and tmr_registers(2)(379)) or                                                       
                            (tmr_registers(0)(379) and tmr_registers(2)(379));                                                         
                                                                                                                                     
        global_tmr_voter(1)(380)  <=    (tmr_registers(0)(380) and tmr_registers(1)(380)) or                                            
                            (tmr_registers(1)(380) and tmr_registers(2)(380)) or                                                       
                            (tmr_registers(0)(380) and tmr_registers(2)(380));                                                         
                                                                                                                                     
        global_tmr_voter(1)(381)  <=    (tmr_registers(0)(381) and tmr_registers(1)(381)) or                                            
                            (tmr_registers(1)(381) and tmr_registers(2)(381)) or                                                       
                            (tmr_registers(0)(381) and tmr_registers(2)(381));                                                         
                                                                                                                                     
        global_tmr_voter(1)(382)  <=    (tmr_registers(0)(382) and tmr_registers(1)(382)) or                                            
                            (tmr_registers(1)(382) and tmr_registers(2)(382)) or                                                       
                            (tmr_registers(0)(382) and tmr_registers(2)(382));                                                         
                                                                                                                                     
        global_tmr_voter(1)(383)  <=    (tmr_registers(0)(383) and tmr_registers(1)(383)) or                                            
                            (tmr_registers(1)(383) and tmr_registers(2)(383)) or                                                       
                            (tmr_registers(0)(383) and tmr_registers(2)(383));                                                         
                                                                                                                                     
        global_tmr_voter(1)(384)  <=    (tmr_registers(0)(384) and tmr_registers(1)(384)) or                                            
                            (tmr_registers(1)(384) and tmr_registers(2)(384)) or                                                       
                            (tmr_registers(0)(384) and tmr_registers(2)(384));                                                         
                                                                                                                                     
        global_tmr_voter(1)(385)  <=    (tmr_registers(0)(385) and tmr_registers(1)(385)) or                                            
                            (tmr_registers(1)(385) and tmr_registers(2)(385)) or                                                       
                            (tmr_registers(0)(385) and tmr_registers(2)(385));                                                         
                                                                                                                                     
        global_tmr_voter(1)(386)  <=    (tmr_registers(0)(386) and tmr_registers(1)(386)) or                                            
                            (tmr_registers(1)(386) and tmr_registers(2)(386)) or                                                       
                            (tmr_registers(0)(386) and tmr_registers(2)(386));                                                         
                                                                                                                                     
        global_tmr_voter(1)(387)  <=    (tmr_registers(0)(387) and tmr_registers(1)(387)) or                                            
                            (tmr_registers(1)(387) and tmr_registers(2)(387)) or                                                       
                            (tmr_registers(0)(387) and tmr_registers(2)(387));                                                         
                                                                                                                                     
        global_tmr_voter(1)(388)  <=    (tmr_registers(0)(388) and tmr_registers(1)(388)) or                                            
                            (tmr_registers(1)(388) and tmr_registers(2)(388)) or                                                       
                            (tmr_registers(0)(388) and tmr_registers(2)(388));                                                         
                                                                                                                                     
        global_tmr_voter(1)(389)  <=    (tmr_registers(0)(389) and tmr_registers(1)(389)) or                                            
                            (tmr_registers(1)(389) and tmr_registers(2)(389)) or                                                       
                            (tmr_registers(0)(389) and tmr_registers(2)(389));                                                         
                                                                                                                                     
        global_tmr_voter(1)(390)  <=    (tmr_registers(0)(390) and tmr_registers(1)(390)) or                                            
                            (tmr_registers(1)(390) and tmr_registers(2)(390)) or                                                       
                            (tmr_registers(0)(390) and tmr_registers(2)(390));                                                         
                                                                                                                                     
        global_tmr_voter(1)(391)  <=    (tmr_registers(0)(391) and tmr_registers(1)(391)) or                                            
                            (tmr_registers(1)(391) and tmr_registers(2)(391)) or                                                       
                            (tmr_registers(0)(391) and tmr_registers(2)(391));                                                         
                                                                                                                                     
        global_tmr_voter(1)(392)  <=    (tmr_registers(0)(392) and tmr_registers(1)(392)) or                                            
                            (tmr_registers(1)(392) and tmr_registers(2)(392)) or                                                       
                            (tmr_registers(0)(392) and tmr_registers(2)(392));                                                         
                                                                                                                                     
        global_tmr_voter(1)(393)  <=    (tmr_registers(0)(393) and tmr_registers(1)(393)) or                                            
                            (tmr_registers(1)(393) and tmr_registers(2)(393)) or                                                       
                            (tmr_registers(0)(393) and tmr_registers(2)(393));                                                         
                                                                                                                                     
        global_tmr_voter(1)(394)  <=    (tmr_registers(0)(394) and tmr_registers(1)(394)) or                                            
                            (tmr_registers(1)(394) and tmr_registers(2)(394)) or                                                       
                            (tmr_registers(0)(394) and tmr_registers(2)(394));                                                         
                                                                                                                                     
        global_tmr_voter(1)(395)  <=    (tmr_registers(0)(395) and tmr_registers(1)(395)) or                                            
                            (tmr_registers(1)(395) and tmr_registers(2)(395)) or                                                       
                            (tmr_registers(0)(395) and tmr_registers(2)(395));                                                         
                                                                                                                                     
        global_tmr_voter(1)(396)  <=    (tmr_registers(0)(396) and tmr_registers(1)(396)) or                                            
                            (tmr_registers(1)(396) and tmr_registers(2)(396)) or                                                       
                            (tmr_registers(0)(396) and tmr_registers(2)(396));                                                         
                                                                                                                                     
        global_tmr_voter(1)(397)  <=    (tmr_registers(0)(397) and tmr_registers(1)(397)) or                                            
                            (tmr_registers(1)(397) and tmr_registers(2)(397)) or                                                       
                            (tmr_registers(0)(397) and tmr_registers(2)(397));                                                         
                                                                                                                                     
        global_tmr_voter(1)(398)  <=    (tmr_registers(0)(398) and tmr_registers(1)(398)) or                                            
                            (tmr_registers(1)(398) and tmr_registers(2)(398)) or                                                       
                            (tmr_registers(0)(398) and tmr_registers(2)(398));                                                         
                                                                                                                                     
        global_tmr_voter(1)(399)  <=    (tmr_registers(0)(399) and tmr_registers(1)(399)) or                                            
                            (tmr_registers(1)(399) and tmr_registers(2)(399)) or                                                       
                            (tmr_registers(0)(399) and tmr_registers(2)(399));                                                         
                                                                                                                                     
        global_tmr_voter(1)(400)  <=    (tmr_registers(0)(400) and tmr_registers(1)(400)) or                                            
                            (tmr_registers(1)(400) and tmr_registers(2)(400)) or                                                       
                            (tmr_registers(0)(400) and tmr_registers(2)(400));                                                         
                                                                                                                                     
        global_tmr_voter(1)(401)  <=    (tmr_registers(0)(401) and tmr_registers(1)(401)) or                                            
                            (tmr_registers(1)(401) and tmr_registers(2)(401)) or                                                       
                            (tmr_registers(0)(401) and tmr_registers(2)(401));                                                         
                                                                                                                                     
        global_tmr_voter(1)(402)  <=    (tmr_registers(0)(402) and tmr_registers(1)(402)) or                                            
                            (tmr_registers(1)(402) and tmr_registers(2)(402)) or                                                       
                            (tmr_registers(0)(402) and tmr_registers(2)(402));                                                         
                                                                                                                                     
        global_tmr_voter(1)(403)  <=    (tmr_registers(0)(403) and tmr_registers(1)(403)) or                                            
                            (tmr_registers(1)(403) and tmr_registers(2)(403)) or                                                       
                            (tmr_registers(0)(403) and tmr_registers(2)(403));                                                         
                                                                                                                                     
        global_tmr_voter(1)(404)  <=    (tmr_registers(0)(404) and tmr_registers(1)(404)) or                                            
                            (tmr_registers(1)(404) and tmr_registers(2)(404)) or                                                       
                            (tmr_registers(0)(404) and tmr_registers(2)(404));                                                         
                                                                                                                                     
        global_tmr_voter(1)(405)  <=    (tmr_registers(0)(405) and tmr_registers(1)(405)) or                                            
                            (tmr_registers(1)(405) and tmr_registers(2)(405)) or                                                       
                            (tmr_registers(0)(405) and tmr_registers(2)(405));                                                         
                                                                                                                                     
        global_tmr_voter(1)(406)  <=    (tmr_registers(0)(406) and tmr_registers(1)(406)) or                                            
                            (tmr_registers(1)(406) and tmr_registers(2)(406)) or                                                       
                            (tmr_registers(0)(406) and tmr_registers(2)(406));                                                         
                                                                                                                                     
        global_tmr_voter(1)(407)  <=    (tmr_registers(0)(407) and tmr_registers(1)(407)) or                                            
                            (tmr_registers(1)(407) and tmr_registers(2)(407)) or                                                       
                            (tmr_registers(0)(407) and tmr_registers(2)(407));                                                         
                                                                                                                                     
        global_tmr_voter(1)(408)  <=    (tmr_registers(0)(408) and tmr_registers(1)(408)) or                                            
                            (tmr_registers(1)(408) and tmr_registers(2)(408)) or                                                       
                            (tmr_registers(0)(408) and tmr_registers(2)(408));                                                         
                                                                                                                                     
        global_tmr_voter(1)(409)  <=    (tmr_registers(0)(409) and tmr_registers(1)(409)) or                                            
                            (tmr_registers(1)(409) and tmr_registers(2)(409)) or                                                       
                            (tmr_registers(0)(409) and tmr_registers(2)(409));                                                         
                                                                                                                                     
        global_tmr_voter(1)(410)  <=    (tmr_registers(0)(410) and tmr_registers(1)(410)) or                                            
                            (tmr_registers(1)(410) and tmr_registers(2)(410)) or                                                       
                            (tmr_registers(0)(410) and tmr_registers(2)(410));                                                         
                                                                                                                                     
        global_tmr_voter(1)(411)  <=    (tmr_registers(0)(411) and tmr_registers(1)(411)) or                                            
                            (tmr_registers(1)(411) and tmr_registers(2)(411)) or                                                       
                            (tmr_registers(0)(411) and tmr_registers(2)(411));                                                         
                                                                                                                                     
        global_tmr_voter(1)(412)  <=    (tmr_registers(0)(412) and tmr_registers(1)(412)) or                                            
                            (tmr_registers(1)(412) and tmr_registers(2)(412)) or                                                       
                            (tmr_registers(0)(412) and tmr_registers(2)(412));                                                         
                                                                                                                                     
        global_tmr_voter(1)(413)  <=    (tmr_registers(0)(413) and tmr_registers(1)(413)) or                                            
                            (tmr_registers(1)(413) and tmr_registers(2)(413)) or                                                       
                            (tmr_registers(0)(413) and tmr_registers(2)(413));                                                         
                                                                                                                                     
        global_tmr_voter(1)(414)  <=    (tmr_registers(0)(414) and tmr_registers(1)(414)) or                                            
                            (tmr_registers(1)(414) and tmr_registers(2)(414)) or                                                       
                            (tmr_registers(0)(414) and tmr_registers(2)(414));                                                         
                                                                                                                                     
        global_tmr_voter(1)(415)  <=    (tmr_registers(0)(415) and tmr_registers(1)(415)) or                                            
                            (tmr_registers(1)(415) and tmr_registers(2)(415)) or                                                       
                            (tmr_registers(0)(415) and tmr_registers(2)(415));                                                         
                                                                                                                                     
        global_tmr_voter(1)(416)  <=    (tmr_registers(0)(416) and tmr_registers(1)(416)) or                                            
                            (tmr_registers(1)(416) and tmr_registers(2)(416)) or                                                       
                            (tmr_registers(0)(416) and tmr_registers(2)(416));                                                         
                                                                                                                                     
        global_tmr_voter(1)(417)  <=    (tmr_registers(0)(417) and tmr_registers(1)(417)) or                                            
                            (tmr_registers(1)(417) and tmr_registers(2)(417)) or                                                       
                            (tmr_registers(0)(417) and tmr_registers(2)(417));                                                         
                                                                                                                                     
        global_tmr_voter(1)(418)  <=    (tmr_registers(0)(418) and tmr_registers(1)(418)) or                                            
                            (tmr_registers(1)(418) and tmr_registers(2)(418)) or                                                       
                            (tmr_registers(0)(418) and tmr_registers(2)(418));                                                         
                                                                                                                                     
        global_tmr_voter(1)(419)  <=    (tmr_registers(0)(419) and tmr_registers(1)(419)) or                                            
                            (tmr_registers(1)(419) and tmr_registers(2)(419)) or                                                       
                            (tmr_registers(0)(419) and tmr_registers(2)(419));                                                         
                                                                                                                                     
        global_tmr_voter(1)(420)  <=    (tmr_registers(0)(420) and tmr_registers(1)(420)) or                                            
                            (tmr_registers(1)(420) and tmr_registers(2)(420)) or                                                       
                            (tmr_registers(0)(420) and tmr_registers(2)(420));                                                         
                                                                                                                                     
        global_tmr_voter(1)(421)  <=    (tmr_registers(0)(421) and tmr_registers(1)(421)) or                                            
                            (tmr_registers(1)(421) and tmr_registers(2)(421)) or                                                       
                            (tmr_registers(0)(421) and tmr_registers(2)(421));                                                         
                                                                                                                                     
        global_tmr_voter(1)(422)  <=    (tmr_registers(0)(422) and tmr_registers(1)(422)) or                                            
                            (tmr_registers(1)(422) and tmr_registers(2)(422)) or                                                       
                            (tmr_registers(0)(422) and tmr_registers(2)(422));                                                         
                                                                                                                                     
        global_tmr_voter(1)(423)  <=    (tmr_registers(0)(423) and tmr_registers(1)(423)) or                                            
                            (tmr_registers(1)(423) and tmr_registers(2)(423)) or                                                       
                            (tmr_registers(0)(423) and tmr_registers(2)(423));                                                         
                                                                                                                                     
        global_tmr_voter(1)(424)  <=    (tmr_registers(0)(424) and tmr_registers(1)(424)) or                                            
                            (tmr_registers(1)(424) and tmr_registers(2)(424)) or                                                       
                            (tmr_registers(0)(424) and tmr_registers(2)(424));                                                         
                                                                                                                                     
        global_tmr_voter(1)(425)  <=    (tmr_registers(0)(425) and tmr_registers(1)(425)) or                                            
                            (tmr_registers(1)(425) and tmr_registers(2)(425)) or                                                       
                            (tmr_registers(0)(425) and tmr_registers(2)(425));                                                         
                                                                                                                                     
        global_tmr_voter(1)(426)  <=    (tmr_registers(0)(426) and tmr_registers(1)(426)) or                                            
                            (tmr_registers(1)(426) and tmr_registers(2)(426)) or                                                       
                            (tmr_registers(0)(426) and tmr_registers(2)(426));                                                         
                                                                                                                                     
        global_tmr_voter(1)(427)  <=    (tmr_registers(0)(427) and tmr_registers(1)(427)) or                                            
                            (tmr_registers(1)(427) and tmr_registers(2)(427)) or                                                       
                            (tmr_registers(0)(427) and tmr_registers(2)(427));                                                         
                                                                                                                                     
        global_tmr_voter(1)(428)  <=    (tmr_registers(0)(428) and tmr_registers(1)(428)) or                                            
                            (tmr_registers(1)(428) and tmr_registers(2)(428)) or                                                       
                            (tmr_registers(0)(428) and tmr_registers(2)(428));                                                         
                                                                                                                                     
        global_tmr_voter(1)(429)  <=    (tmr_registers(0)(429) and tmr_registers(1)(429)) or                                            
                            (tmr_registers(1)(429) and tmr_registers(2)(429)) or                                                       
                            (tmr_registers(0)(429) and tmr_registers(2)(429));                                                         
                                                                                                                                     
        global_tmr_voter(1)(430)  <=    (tmr_registers(0)(430) and tmr_registers(1)(430)) or                                            
                            (tmr_registers(1)(430) and tmr_registers(2)(430)) or                                                       
                            (tmr_registers(0)(430) and tmr_registers(2)(430));                                                         
                                                                                                                                     
        global_tmr_voter(1)(431)  <=    (tmr_registers(0)(431) and tmr_registers(1)(431)) or                                            
                            (tmr_registers(1)(431) and tmr_registers(2)(431)) or                                                       
                            (tmr_registers(0)(431) and tmr_registers(2)(431));                                                         
                                                                                                                                     
        global_tmr_voter(1)(432)  <=    (tmr_registers(0)(432) and tmr_registers(1)(432)) or                                            
                            (tmr_registers(1)(432) and tmr_registers(2)(432)) or                                                       
                            (tmr_registers(0)(432) and tmr_registers(2)(432));                                                         
                                                                                                                                     
        global_tmr_voter(1)(433)  <=    (tmr_registers(0)(433) and tmr_registers(1)(433)) or                                            
                            (tmr_registers(1)(433) and tmr_registers(2)(433)) or                                                       
                            (tmr_registers(0)(433) and tmr_registers(2)(433));                                                         
                                                                                                                                     
        global_tmr_voter(1)(434)  <=    (tmr_registers(0)(434) and tmr_registers(1)(434)) or                                            
                            (tmr_registers(1)(434) and tmr_registers(2)(434)) or                                                       
                            (tmr_registers(0)(434) and tmr_registers(2)(434));                                                         
                                                                                                                                     
        global_tmr_voter(1)(435)  <=    (tmr_registers(0)(435) and tmr_registers(1)(435)) or                                            
                            (tmr_registers(1)(435) and tmr_registers(2)(435)) or                                                       
                            (tmr_registers(0)(435) and tmr_registers(2)(435));                                                         
                                                                                                                                     
        global_tmr_voter(1)(436)  <=    (tmr_registers(0)(436) and tmr_registers(1)(436)) or                                            
                            (tmr_registers(1)(436) and tmr_registers(2)(436)) or                                                       
                            (tmr_registers(0)(436) and tmr_registers(2)(436));                                                         
                                                                                                                                     
        global_tmr_voter(1)(437)  <=    (tmr_registers(0)(437) and tmr_registers(1)(437)) or                                            
                            (tmr_registers(1)(437) and tmr_registers(2)(437)) or                                                       
                            (tmr_registers(0)(437) and tmr_registers(2)(437));                                                         
                                                                                                                                     
        global_tmr_voter(1)(438)  <=    (tmr_registers(0)(438) and tmr_registers(1)(438)) or                                            
                            (tmr_registers(1)(438) and tmr_registers(2)(438)) or                                                       
                            (tmr_registers(0)(438) and tmr_registers(2)(438));                                                         
                                                                                                                                     
        global_tmr_voter(1)(439)  <=    (tmr_registers(0)(439) and tmr_registers(1)(439)) or                                            
                            (tmr_registers(1)(439) and tmr_registers(2)(439)) or                                                       
                            (tmr_registers(0)(439) and tmr_registers(2)(439));                                                         
                                                                                                                                     
        global_tmr_voter(1)(440)  <=    (tmr_registers(0)(440) and tmr_registers(1)(440)) or                                            
                            (tmr_registers(1)(440) and tmr_registers(2)(440)) or                                                       
                            (tmr_registers(0)(440) and tmr_registers(2)(440));                                                         
                                                                                                                                     
        global_tmr_voter(1)(441)  <=    (tmr_registers(0)(441) and tmr_registers(1)(441)) or                                            
                            (tmr_registers(1)(441) and tmr_registers(2)(441)) or                                                       
                            (tmr_registers(0)(441) and tmr_registers(2)(441));                                                         
                                                                                                                                     
        global_tmr_voter(1)(442)  <=    (tmr_registers(0)(442) and tmr_registers(1)(442)) or                                            
                            (tmr_registers(1)(442) and tmr_registers(2)(442)) or                                                       
                            (tmr_registers(0)(442) and tmr_registers(2)(442));                                                         
                                                                                                                                     
        global_tmr_voter(1)(443)  <=    (tmr_registers(0)(443) and tmr_registers(1)(443)) or                                            
                            (tmr_registers(1)(443) and tmr_registers(2)(443)) or                                                       
                            (tmr_registers(0)(443) and tmr_registers(2)(443));                                                         
                                                                                                                                     
        global_tmr_voter(1)(444)  <=    (tmr_registers(0)(444) and tmr_registers(1)(444)) or                                            
                            (tmr_registers(1)(444) and tmr_registers(2)(444)) or                                                       
                            (tmr_registers(0)(444) and tmr_registers(2)(444));                                                         
                                                                                                                                     
        global_tmr_voter(1)(445)  <=    (tmr_registers(0)(445) and tmr_registers(1)(445)) or                                            
                            (tmr_registers(1)(445) and tmr_registers(2)(445)) or                                                       
                            (tmr_registers(0)(445) and tmr_registers(2)(445));                                                         
                                                                                                                                     
        global_tmr_voter(1)(446)  <=    (tmr_registers(0)(446) and tmr_registers(1)(446)) or                                            
                            (tmr_registers(1)(446) and tmr_registers(2)(446)) or                                                       
                            (tmr_registers(0)(446) and tmr_registers(2)(446));                                                         
                                                                                                                                     
        global_tmr_voter(1)(447)  <=    (tmr_registers(0)(447) and tmr_registers(1)(447)) or                                            
                            (tmr_registers(1)(447) and tmr_registers(2)(447)) or                                                       
                            (tmr_registers(0)(447) and tmr_registers(2)(447));                                                         
                                                                                                                                     
        global_tmr_voter(1)(448)  <=    (tmr_registers(0)(448) and tmr_registers(1)(448)) or                                            
                            (tmr_registers(1)(448) and tmr_registers(2)(448)) or                                                       
                            (tmr_registers(0)(448) and tmr_registers(2)(448));                                                         
                                                                                                                                     
        global_tmr_voter(1)(449)  <=    (tmr_registers(0)(449) and tmr_registers(1)(449)) or                                            
                            (tmr_registers(1)(449) and tmr_registers(2)(449)) or                                                       
                            (tmr_registers(0)(449) and tmr_registers(2)(449));                                                         
                                                                                                                                     
        global_tmr_voter(1)(450)  <=    (tmr_registers(0)(450) and tmr_registers(1)(450)) or                                            
                            (tmr_registers(1)(450) and tmr_registers(2)(450)) or                                                       
                            (tmr_registers(0)(450) and tmr_registers(2)(450));                                                         
                                                                                                                                     
        global_tmr_voter(1)(451)  <=    (tmr_registers(0)(451) and tmr_registers(1)(451)) or                                            
                            (tmr_registers(1)(451) and tmr_registers(2)(451)) or                                                       
                            (tmr_registers(0)(451) and tmr_registers(2)(451));                                                         
                                                                                                                                     
        global_tmr_voter(1)(452)  <=    (tmr_registers(0)(452) and tmr_registers(1)(452)) or                                            
                            (tmr_registers(1)(452) and tmr_registers(2)(452)) or                                                       
                            (tmr_registers(0)(452) and tmr_registers(2)(452));                                                         
                                                                                                                                     
        global_tmr_voter(1)(453)  <=    (tmr_registers(0)(453) and tmr_registers(1)(453)) or                                            
                            (tmr_registers(1)(453) and tmr_registers(2)(453)) or                                                       
                            (tmr_registers(0)(453) and tmr_registers(2)(453));                                                         
                                                                                                                                     
        global_tmr_voter(1)(454)  <=    (tmr_registers(0)(454) and tmr_registers(1)(454)) or                                            
                            (tmr_registers(1)(454) and tmr_registers(2)(454)) or                                                       
                            (tmr_registers(0)(454) and tmr_registers(2)(454));                                                         
                                                                                                                                     
        global_tmr_voter(1)(455)  <=    (tmr_registers(0)(455) and tmr_registers(1)(455)) or                                            
                            (tmr_registers(1)(455) and tmr_registers(2)(455)) or                                                       
                            (tmr_registers(0)(455) and tmr_registers(2)(455));                                                         
                                                                                                                                     
        global_tmr_voter(1)(456)  <=    (tmr_registers(0)(456) and tmr_registers(1)(456)) or                                            
                            (tmr_registers(1)(456) and tmr_registers(2)(456)) or                                                       
                            (tmr_registers(0)(456) and tmr_registers(2)(456));                                                         
                                                                                                                                     
        global_tmr_voter(1)(457)  <=    (tmr_registers(0)(457) and tmr_registers(1)(457)) or                                            
                            (tmr_registers(1)(457) and tmr_registers(2)(457)) or                                                       
                            (tmr_registers(0)(457) and tmr_registers(2)(457));                                                         
                                                                                                                                     
        global_tmr_voter(1)(458)  <=    (tmr_registers(0)(458) and tmr_registers(1)(458)) or                                            
                            (tmr_registers(1)(458) and tmr_registers(2)(458)) or                                                       
                            (tmr_registers(0)(458) and tmr_registers(2)(458));                                                         
                                                                                                                                     
        global_tmr_voter(1)(459)  <=    (tmr_registers(0)(459) and tmr_registers(1)(459)) or                                            
                            (tmr_registers(1)(459) and tmr_registers(2)(459)) or                                                       
                            (tmr_registers(0)(459) and tmr_registers(2)(459));                                                         
                                                                                                                                     
        global_tmr_voter(1)(460)  <=    (tmr_registers(0)(460) and tmr_registers(1)(460)) or                                            
                            (tmr_registers(1)(460) and tmr_registers(2)(460)) or                                                       
                            (tmr_registers(0)(460) and tmr_registers(2)(460));                                                         
                                                                                                                                     
        global_tmr_voter(1)(461)  <=    (tmr_registers(0)(461) and tmr_registers(1)(461)) or                                            
                            (tmr_registers(1)(461) and tmr_registers(2)(461)) or                                                       
                            (tmr_registers(0)(461) and tmr_registers(2)(461));                                                         
                                                                                                                                     
        global_tmr_voter(1)(462)  <=    (tmr_registers(0)(462) and tmr_registers(1)(462)) or                                            
                            (tmr_registers(1)(462) and tmr_registers(2)(462)) or                                                       
                            (tmr_registers(0)(462) and tmr_registers(2)(462));                                                         
                                                                                                                                     
        global_tmr_voter(1)(463)  <=    (tmr_registers(0)(463) and tmr_registers(1)(463)) or                                            
                            (tmr_registers(1)(463) and tmr_registers(2)(463)) or                                                       
                            (tmr_registers(0)(463) and tmr_registers(2)(463));                                                         
                                                                                                                                     
        global_tmr_voter(1)(464)  <=    (tmr_registers(0)(464) and tmr_registers(1)(464)) or                                            
                            (tmr_registers(1)(464) and tmr_registers(2)(464)) or                                                       
                            (tmr_registers(0)(464) and tmr_registers(2)(464));                                                         
                                                                                                                                     
        global_tmr_voter(1)(465)  <=    (tmr_registers(0)(465) and tmr_registers(1)(465)) or                                            
                            (tmr_registers(1)(465) and tmr_registers(2)(465)) or                                                       
                            (tmr_registers(0)(465) and tmr_registers(2)(465));                                                         
                                                                                                                                     
        global_tmr_voter(1)(466)  <=    (tmr_registers(0)(466) and tmr_registers(1)(466)) or                                            
                            (tmr_registers(1)(466) and tmr_registers(2)(466)) or                                                       
                            (tmr_registers(0)(466) and tmr_registers(2)(466));                                                         
                                                                                                                                     
        global_tmr_voter(1)(467)  <=    (tmr_registers(0)(467) and tmr_registers(1)(467)) or                                            
                            (tmr_registers(1)(467) and tmr_registers(2)(467)) or                                                       
                            (tmr_registers(0)(467) and tmr_registers(2)(467));                                                         
                                                                                                                                     
        global_tmr_voter(1)(468)  <=    (tmr_registers(0)(468) and tmr_registers(1)(468)) or                                            
                            (tmr_registers(1)(468) and tmr_registers(2)(468)) or                                                       
                            (tmr_registers(0)(468) and tmr_registers(2)(468));                                                         
                                                                                                                                     
        global_tmr_voter(1)(469)  <=    (tmr_registers(0)(469) and tmr_registers(1)(469)) or                                            
                            (tmr_registers(1)(469) and tmr_registers(2)(469)) or                                                       
                            (tmr_registers(0)(469) and tmr_registers(2)(469));                                                         
                                                                                                                                     
        global_tmr_voter(1)(470)  <=    (tmr_registers(0)(470) and tmr_registers(1)(470)) or                                            
                            (tmr_registers(1)(470) and tmr_registers(2)(470)) or                                                       
                            (tmr_registers(0)(470) and tmr_registers(2)(470));                                                         
                                                                                                                                     
        global_tmr_voter(1)(471)  <=    (tmr_registers(0)(471) and tmr_registers(1)(471)) or                                            
                            (tmr_registers(1)(471) and tmr_registers(2)(471)) or                                                       
                            (tmr_registers(0)(471) and tmr_registers(2)(471));                                                         
                                                                                                                                     
        global_tmr_voter(1)(472)  <=    (tmr_registers(0)(472) and tmr_registers(1)(472)) or                                            
                            (tmr_registers(1)(472) and tmr_registers(2)(472)) or                                                       
                            (tmr_registers(0)(472) and tmr_registers(2)(472));                                                         
                                                                                                                                     
        global_tmr_voter(1)(473)  <=    (tmr_registers(0)(473) and tmr_registers(1)(473)) or                                            
                            (tmr_registers(1)(473) and tmr_registers(2)(473)) or                                                       
                            (tmr_registers(0)(473) and tmr_registers(2)(473));                                                         
                                                                                                                                     
        global_tmr_voter(1)(474)  <=    (tmr_registers(0)(474) and tmr_registers(1)(474)) or                                            
                            (tmr_registers(1)(474) and tmr_registers(2)(474)) or                                                       
                            (tmr_registers(0)(474) and tmr_registers(2)(474));                                                         
                                                                                                                                     
        global_tmr_voter(1)(475)  <=    (tmr_registers(0)(475) and tmr_registers(1)(475)) or                                            
                            (tmr_registers(1)(475) and tmr_registers(2)(475)) or                                                       
                            (tmr_registers(0)(475) and tmr_registers(2)(475));                                                         
                                                                                                                                     
        global_tmr_voter(1)(476)  <=    (tmr_registers(0)(476) and tmr_registers(1)(476)) or                                            
                            (tmr_registers(1)(476) and tmr_registers(2)(476)) or                                                       
                            (tmr_registers(0)(476) and tmr_registers(2)(476));                                                         
                                                                                                                                     
        global_tmr_voter(1)(477)  <=    (tmr_registers(0)(477) and tmr_registers(1)(477)) or                                            
                            (tmr_registers(1)(477) and tmr_registers(2)(477)) or                                                       
                            (tmr_registers(0)(477) and tmr_registers(2)(477));                                                         
                                                                                                                                     
        global_tmr_voter(1)(478)  <=    (tmr_registers(0)(478) and tmr_registers(1)(478)) or                                            
                            (tmr_registers(1)(478) and tmr_registers(2)(478)) or                                                       
                            (tmr_registers(0)(478) and tmr_registers(2)(478));                                                         
                                                                                                                                     
        global_tmr_voter(1)(479)  <=    (tmr_registers(0)(479) and tmr_registers(1)(479)) or                                            
                            (tmr_registers(1)(479) and tmr_registers(2)(479)) or                                                       
                            (tmr_registers(0)(479) and tmr_registers(2)(479));                                                         
                                                                                                                                     
        global_tmr_voter(1)(480)  <=    (tmr_registers(0)(480) and tmr_registers(1)(480)) or                                            
                            (tmr_registers(1)(480) and tmr_registers(2)(480)) or                                                       
                            (tmr_registers(0)(480) and tmr_registers(2)(480));                                                         
                                                                                                                                     
        global_tmr_voter(1)(481)  <=    (tmr_registers(0)(481) and tmr_registers(1)(481)) or                                            
                            (tmr_registers(1)(481) and tmr_registers(2)(481)) or                                                       
                            (tmr_registers(0)(481) and tmr_registers(2)(481));                                                         
                                                                                                                                     
        global_tmr_voter(1)(482)  <=    (tmr_registers(0)(482) and tmr_registers(1)(482)) or                                            
                            (tmr_registers(1)(482) and tmr_registers(2)(482)) or                                                       
                            (tmr_registers(0)(482) and tmr_registers(2)(482));                                                         
                                                                                                                                     
        global_tmr_voter(1)(483)  <=    (tmr_registers(0)(483) and tmr_registers(1)(483)) or                                            
                            (tmr_registers(1)(483) and tmr_registers(2)(483)) or                                                       
                            (tmr_registers(0)(483) and tmr_registers(2)(483));                                                         
                                                                                                                                     
        global_tmr_voter(1)(484)  <=    (tmr_registers(0)(484) and tmr_registers(1)(484)) or                                            
                            (tmr_registers(1)(484) and tmr_registers(2)(484)) or                                                       
                            (tmr_registers(0)(484) and tmr_registers(2)(484));                                                         
                                                                                                                                     
        global_tmr_voter(1)(485)  <=    (tmr_registers(0)(485) and tmr_registers(1)(485)) or                                            
                            (tmr_registers(1)(485) and tmr_registers(2)(485)) or                                                       
                            (tmr_registers(0)(485) and tmr_registers(2)(485));                                                         
                                                                                                                                     
        global_tmr_voter(1)(486)  <=    (tmr_registers(0)(486) and tmr_registers(1)(486)) or                                            
                            (tmr_registers(1)(486) and tmr_registers(2)(486)) or                                                       
                            (tmr_registers(0)(486) and tmr_registers(2)(486));                                                         
                                                                                                                                     
        global_tmr_voter(1)(487)  <=    (tmr_registers(0)(487) and tmr_registers(1)(487)) or                                            
                            (tmr_registers(1)(487) and tmr_registers(2)(487)) or                                                       
                            (tmr_registers(0)(487) and tmr_registers(2)(487));                                                         
                                                                                                                                     
        global_tmr_voter(1)(488)  <=    (tmr_registers(0)(488) and tmr_registers(1)(488)) or                                            
                            (tmr_registers(1)(488) and tmr_registers(2)(488)) or                                                       
                            (tmr_registers(0)(488) and tmr_registers(2)(488));                                                         
                                                                                                                                     
        global_tmr_voter(1)(489)  <=    (tmr_registers(0)(489) and tmr_registers(1)(489)) or                                            
                            (tmr_registers(1)(489) and tmr_registers(2)(489)) or                                                       
                            (tmr_registers(0)(489) and tmr_registers(2)(489));                                                         
                                                                                                                                     
        global_tmr_voter(1)(490)  <=    (tmr_registers(0)(490) and tmr_registers(1)(490)) or                                            
                            (tmr_registers(1)(490) and tmr_registers(2)(490)) or                                                       
                            (tmr_registers(0)(490) and tmr_registers(2)(490));                                                         
                                                                                                                                     
        global_tmr_voter(1)(491)  <=    (tmr_registers(0)(491) and tmr_registers(1)(491)) or                                            
                            (tmr_registers(1)(491) and tmr_registers(2)(491)) or                                                       
                            (tmr_registers(0)(491) and tmr_registers(2)(491));                                                         
                                                                                                                                     
        global_tmr_voter(1)(492)  <=    (tmr_registers(0)(492) and tmr_registers(1)(492)) or                                            
                            (tmr_registers(1)(492) and tmr_registers(2)(492)) or                                                       
                            (tmr_registers(0)(492) and tmr_registers(2)(492));                                                         
                                                                                                                                     
        global_tmr_voter(1)(493)  <=    (tmr_registers(0)(493) and tmr_registers(1)(493)) or                                            
                            (tmr_registers(1)(493) and tmr_registers(2)(493)) or                                                       
                            (tmr_registers(0)(493) and tmr_registers(2)(493));                                                         
                                                                                                                                     
        global_tmr_voter(1)(494)  <=    (tmr_registers(0)(494) and tmr_registers(1)(494)) or                                            
                            (tmr_registers(1)(494) and tmr_registers(2)(494)) or                                                       
                            (tmr_registers(0)(494) and tmr_registers(2)(494));                                                         
                                                                                                                                     
        global_tmr_voter(1)(495)  <=    (tmr_registers(0)(495) and tmr_registers(1)(495)) or                                            
                            (tmr_registers(1)(495) and tmr_registers(2)(495)) or                                                       
                            (tmr_registers(0)(495) and tmr_registers(2)(495));                                                         
                                                                                                                                     
        global_tmr_voter(1)(496)  <=    (tmr_registers(0)(496) and tmr_registers(1)(496)) or                                            
                            (tmr_registers(1)(496) and tmr_registers(2)(496)) or                                                       
                            (tmr_registers(0)(496) and tmr_registers(2)(496));                                                         
                                                                                                                                     
        global_tmr_voter(1)(497)  <=    (tmr_registers(0)(497) and tmr_registers(1)(497)) or                                            
                            (tmr_registers(1)(497) and tmr_registers(2)(497)) or                                                       
                            (tmr_registers(0)(497) and tmr_registers(2)(497));                                                         
                                                                                                                                     
        global_tmr_voter(1)(498)  <=    (tmr_registers(0)(498) and tmr_registers(1)(498)) or                                            
                            (tmr_registers(1)(498) and tmr_registers(2)(498)) or                                                       
                            (tmr_registers(0)(498) and tmr_registers(2)(498));                                                         
                                                                                                                                     
        global_tmr_voter(1)(499)  <=    (tmr_registers(0)(499) and tmr_registers(1)(499)) or                                            
                            (tmr_registers(1)(499) and tmr_registers(2)(499)) or                                                       
                            (tmr_registers(0)(499) and tmr_registers(2)(499));                                                         
                                                                                                                                     
        global_tmr_voter(1)(500)  <=    (tmr_registers(0)(500) and tmr_registers(1)(500)) or                                            
                            (tmr_registers(1)(500) and tmr_registers(2)(500)) or                                                       
                            (tmr_registers(0)(500) and tmr_registers(2)(500));                                                         
                                                                                                                                     
        global_tmr_voter(1)(501)  <=    (tmr_registers(0)(501) and tmr_registers(1)(501)) or                                            
                            (tmr_registers(1)(501) and tmr_registers(2)(501)) or                                                       
                            (tmr_registers(0)(501) and tmr_registers(2)(501));                                                         
                                                                                                                                     
        global_tmr_voter(1)(502)  <=    (tmr_registers(0)(502) and tmr_registers(1)(502)) or                                            
                            (tmr_registers(1)(502) and tmr_registers(2)(502)) or                                                       
                            (tmr_registers(0)(502) and tmr_registers(2)(502));                                                         
                                                                                                                                     
        global_tmr_voter(1)(503)  <=    (tmr_registers(0)(503) and tmr_registers(1)(503)) or                                            
                            (tmr_registers(1)(503) and tmr_registers(2)(503)) or                                                       
                            (tmr_registers(0)(503) and tmr_registers(2)(503));                                                         
                                                                                                                                     
        global_tmr_voter(1)(504)  <=    (tmr_registers(0)(504) and tmr_registers(1)(504)) or                                            
                            (tmr_registers(1)(504) and tmr_registers(2)(504)) or                                                       
                            (tmr_registers(0)(504) and tmr_registers(2)(504));                                                         
                                                                                                                                     
        global_tmr_voter(1)(505)  <=    (tmr_registers(0)(505) and tmr_registers(1)(505)) or                                            
                            (tmr_registers(1)(505) and tmr_registers(2)(505)) or                                                       
                            (tmr_registers(0)(505) and tmr_registers(2)(505));                                                         
                                                                                                                                     
        global_tmr_voter(1)(506)  <=    (tmr_registers(0)(506) and tmr_registers(1)(506)) or                                            
                            (tmr_registers(1)(506) and tmr_registers(2)(506)) or                                                       
                            (tmr_registers(0)(506) and tmr_registers(2)(506));                                                         
                                                                                                                                     
        global_tmr_voter(1)(507)  <=    (tmr_registers(0)(507) and tmr_registers(1)(507)) or                                            
                            (tmr_registers(1)(507) and tmr_registers(2)(507)) or                                                       
                            (tmr_registers(0)(507) and tmr_registers(2)(507));                                                         
                                                                                                                                     
        global_tmr_voter(1)(508)  <=    (tmr_registers(0)(508) and tmr_registers(1)(508)) or                                            
                            (tmr_registers(1)(508) and tmr_registers(2)(508)) or                                                       
                            (tmr_registers(0)(508) and tmr_registers(2)(508));                                                         
                                                                                                                                     
        global_tmr_voter(1)(509)  <=    (tmr_registers(0)(509) and tmr_registers(1)(509)) or                                            
                            (tmr_registers(1)(509) and tmr_registers(2)(509)) or                                                       
                            (tmr_registers(0)(509) and tmr_registers(2)(509));                                                         
                                                                                                                                     
        global_tmr_voter(1)(510)  <=    (tmr_registers(0)(510) and tmr_registers(1)(510)) or                                            
                            (tmr_registers(1)(510) and tmr_registers(2)(510)) or                                                       
                            (tmr_registers(0)(510) and tmr_registers(2)(510));                                                         
                                                                                                                                     
        global_tmr_voter(1)(511)  <=    (tmr_registers(0)(511) and tmr_registers(1)(511)) or                                            
                            (tmr_registers(1)(511) and tmr_registers(2)(511)) or                                                       
                            (tmr_registers(0)(511) and tmr_registers(2)(511));                                                         
                                                                                                                                     
        global_tmr_voter(1)(512)  <=    (tmr_registers(0)(512) and tmr_registers(1)(512)) or                                            
                            (tmr_registers(1)(512) and tmr_registers(2)(512)) or                                                       
                            (tmr_registers(0)(512) and tmr_registers(2)(512));                                                         
                                                                                                                                     
        global_tmr_voter(1)(513)  <=    (tmr_registers(0)(513) and tmr_registers(1)(513)) or                                            
                            (tmr_registers(1)(513) and tmr_registers(2)(513)) or                                                       
                            (tmr_registers(0)(513) and tmr_registers(2)(513));                                                         
                                                                                                                                     
        global_tmr_voter(1)(514)  <=    (tmr_registers(0)(514) and tmr_registers(1)(514)) or                                            
                            (tmr_registers(1)(514) and tmr_registers(2)(514)) or                                                       
                            (tmr_registers(0)(514) and tmr_registers(2)(514));                                                         
                                                                                                                                     
        global_tmr_voter(1)(515)  <=    (tmr_registers(0)(515) and tmr_registers(1)(515)) or                                            
                            (tmr_registers(1)(515) and tmr_registers(2)(515)) or                                                       
                            (tmr_registers(0)(515) and tmr_registers(2)(515));                                                         
                                                                                                                                     
        global_tmr_voter(1)(516)  <=    (tmr_registers(0)(516) and tmr_registers(1)(516)) or                                            
                            (tmr_registers(1)(516) and tmr_registers(2)(516)) or                                                       
                            (tmr_registers(0)(516) and tmr_registers(2)(516));                                                         
                                                                                                                                     
        global_tmr_voter(1)(517)  <=    (tmr_registers(0)(517) and tmr_registers(1)(517)) or                                            
                            (tmr_registers(1)(517) and tmr_registers(2)(517)) or                                                       
                            (tmr_registers(0)(517) and tmr_registers(2)(517));                                                         
                                                                                                                                     
        global_tmr_voter(1)(518)  <=    (tmr_registers(0)(518) and tmr_registers(1)(518)) or                                            
                            (tmr_registers(1)(518) and tmr_registers(2)(518)) or                                                       
                            (tmr_registers(0)(518) and tmr_registers(2)(518));                                                         
                                                                                                                                     
        global_tmr_voter(1)(519)  <=    (tmr_registers(0)(519) and tmr_registers(1)(519)) or                                            
                            (tmr_registers(1)(519) and tmr_registers(2)(519)) or                                                       
                            (tmr_registers(0)(519) and tmr_registers(2)(519));                                                         
                                                                                                                                     
        global_tmr_voter(1)(520)  <=    (tmr_registers(0)(520) and tmr_registers(1)(520)) or                                            
                            (tmr_registers(1)(520) and tmr_registers(2)(520)) or                                                       
                            (tmr_registers(0)(520) and tmr_registers(2)(520));                                                         
                                                                                                                                     
        global_tmr_voter(1)(521)  <=    (tmr_registers(0)(521) and tmr_registers(1)(521)) or                                            
                            (tmr_registers(1)(521) and tmr_registers(2)(521)) or                                                       
                            (tmr_registers(0)(521) and tmr_registers(2)(521));                                                         
                                                                                                                                     
        global_tmr_voter(1)(522)  <=    (tmr_registers(0)(522) and tmr_registers(1)(522)) or                                            
                            (tmr_registers(1)(522) and tmr_registers(2)(522)) or                                                       
                            (tmr_registers(0)(522) and tmr_registers(2)(522));                                                         
                                                                                                                                     
        global_tmr_voter(1)(523)  <=    (tmr_registers(0)(523) and tmr_registers(1)(523)) or                                            
                            (tmr_registers(1)(523) and tmr_registers(2)(523)) or                                                       
                            (tmr_registers(0)(523) and tmr_registers(2)(523));                                                         
                                                                                                                                     
        global_tmr_voter(1)(524)  <=    (tmr_registers(0)(524) and tmr_registers(1)(524)) or                                            
                            (tmr_registers(1)(524) and tmr_registers(2)(524)) or                                                       
                            (tmr_registers(0)(524) and tmr_registers(2)(524));                                                         
                                                                                                                                     
        global_tmr_voter(1)(525)  <=    (tmr_registers(0)(525) and tmr_registers(1)(525)) or                                            
                            (tmr_registers(1)(525) and tmr_registers(2)(525)) or                                                       
                            (tmr_registers(0)(525) and tmr_registers(2)(525));                                                         
                                                                                                                                     
        global_tmr_voter(1)(526)  <=    (tmr_registers(0)(526) and tmr_registers(1)(526)) or                                            
                            (tmr_registers(1)(526) and tmr_registers(2)(526)) or                                                       
                            (tmr_registers(0)(526) and tmr_registers(2)(526));                                                         
                                                                                                                                     
        global_tmr_voter(1)(527)  <=    (tmr_registers(0)(527) and tmr_registers(1)(527)) or                                            
                            (tmr_registers(1)(527) and tmr_registers(2)(527)) or                                                       
                            (tmr_registers(0)(527) and tmr_registers(2)(527));                                                         
                                                                                                                                     
        global_tmr_voter(1)(528)  <=    (tmr_registers(0)(528) and tmr_registers(1)(528)) or                                            
                            (tmr_registers(1)(528) and tmr_registers(2)(528)) or                                                       
                            (tmr_registers(0)(528) and tmr_registers(2)(528));                                                         
                                                                                                                                     
        global_tmr_voter(1)(529)  <=    (tmr_registers(0)(529) and tmr_registers(1)(529)) or                                            
                            (tmr_registers(1)(529) and tmr_registers(2)(529)) or                                                       
                            (tmr_registers(0)(529) and tmr_registers(2)(529));                                                         
                                                                                                                                     
        global_tmr_voter(1)(530)  <=    (tmr_registers(0)(530) and tmr_registers(1)(530)) or                                            
                            (tmr_registers(1)(530) and tmr_registers(2)(530)) or                                                       
                            (tmr_registers(0)(530) and tmr_registers(2)(530));                                                         
                                                                                                                                     
        global_tmr_voter(1)(531)  <=    (tmr_registers(0)(531) and tmr_registers(1)(531)) or                                            
                            (tmr_registers(1)(531) and tmr_registers(2)(531)) or                                                       
                            (tmr_registers(0)(531) and tmr_registers(2)(531));                                                         
                                                                                                                                     
        global_tmr_voter(1)(532)  <=    (tmr_registers(0)(532) and tmr_registers(1)(532)) or                                            
                            (tmr_registers(1)(532) and tmr_registers(2)(532)) or                                                       
                            (tmr_registers(0)(532) and tmr_registers(2)(532));                                                         
                                                                                                                                     
        global_tmr_voter(1)(533)  <=    (tmr_registers(0)(533) and tmr_registers(1)(533)) or                                            
                            (tmr_registers(1)(533) and tmr_registers(2)(533)) or                                                       
                            (tmr_registers(0)(533) and tmr_registers(2)(533));                                                         
                                                                                                                                     
        global_tmr_voter(1)(534)  <=    (tmr_registers(0)(534) and tmr_registers(1)(534)) or                                            
                            (tmr_registers(1)(534) and tmr_registers(2)(534)) or                                                       
                            (tmr_registers(0)(534) and tmr_registers(2)(534));                                                         
                                                                                                                                     
        global_tmr_voter(1)(535)  <=    (tmr_registers(0)(535) and tmr_registers(1)(535)) or                                            
                            (tmr_registers(1)(535) and tmr_registers(2)(535)) or                                                       
                            (tmr_registers(0)(535) and tmr_registers(2)(535));                                                         
                                                                                                                                     
        global_tmr_voter(1)(536)  <=    (tmr_registers(0)(536) and tmr_registers(1)(536)) or                                            
                            (tmr_registers(1)(536) and tmr_registers(2)(536)) or                                                       
                            (tmr_registers(0)(536) and tmr_registers(2)(536));                                                         
                                                                                                                                     
        global_tmr_voter(1)(537)  <=    (tmr_registers(0)(537) and tmr_registers(1)(537)) or                                            
                            (tmr_registers(1)(537) and tmr_registers(2)(537)) or                                                       
                            (tmr_registers(0)(537) and tmr_registers(2)(537));                                                         
                                                                                                                                     
        global_tmr_voter(1)(538)  <=    (tmr_registers(0)(538) and tmr_registers(1)(538)) or                                            
                            (tmr_registers(1)(538) and tmr_registers(2)(538)) or                                                       
                            (tmr_registers(0)(538) and tmr_registers(2)(538));                                                         
                                                                                                                                     
        global_tmr_voter(1)(539)  <=    (tmr_registers(0)(539) and tmr_registers(1)(539)) or                                            
                            (tmr_registers(1)(539) and tmr_registers(2)(539)) or                                                       
                            (tmr_registers(0)(539) and tmr_registers(2)(539));                                                         
                                                                                                                                     
        global_tmr_voter(1)(540)  <=    (tmr_registers(0)(540) and tmr_registers(1)(540)) or                                            
                            (tmr_registers(1)(540) and tmr_registers(2)(540)) or                                                       
                            (tmr_registers(0)(540) and tmr_registers(2)(540));                                                         
                                                                                                                                     
        global_tmr_voter(1)(541)  <=    (tmr_registers(0)(541) and tmr_registers(1)(541)) or                                            
                            (tmr_registers(1)(541) and tmr_registers(2)(541)) or                                                       
                            (tmr_registers(0)(541) and tmr_registers(2)(541));                                                         
                                                                                                                                     
        global_tmr_voter(1)(542)  <=    (tmr_registers(0)(542) and tmr_registers(1)(542)) or                                            
                            (tmr_registers(1)(542) and tmr_registers(2)(542)) or                                                       
                            (tmr_registers(0)(542) and tmr_registers(2)(542));                                                         
                                                                                                                                     
        global_tmr_voter(1)(543)  <=    (tmr_registers(0)(543) and tmr_registers(1)(543)) or                                            
                            (tmr_registers(1)(543) and tmr_registers(2)(543)) or                                                       
                            (tmr_registers(0)(543) and tmr_registers(2)(543));                                                         
                                                                                                                                     
        global_tmr_voter(1)(544)  <=    (tmr_registers(0)(544) and tmr_registers(1)(544)) or                                            
                            (tmr_registers(1)(544) and tmr_registers(2)(544)) or                                                       
                            (tmr_registers(0)(544) and tmr_registers(2)(544));                                                         
                                                                                                                                     
        global_tmr_voter(1)(545)  <=    (tmr_registers(0)(545) and tmr_registers(1)(545)) or                                            
                            (tmr_registers(1)(545) and tmr_registers(2)(545)) or                                                       
                            (tmr_registers(0)(545) and tmr_registers(2)(545));                                                         
                                                                                                                                     
        global_tmr_voter(1)(546)  <=    (tmr_registers(0)(546) and tmr_registers(1)(546)) or                                            
                            (tmr_registers(1)(546) and tmr_registers(2)(546)) or                                                       
                            (tmr_registers(0)(546) and tmr_registers(2)(546));                                                         
                                                                                                                                     
        global_tmr_voter(1)(547)  <=    (tmr_registers(0)(547) and tmr_registers(1)(547)) or                                            
                            (tmr_registers(1)(547) and tmr_registers(2)(547)) or                                                       
                            (tmr_registers(0)(547) and tmr_registers(2)(547));                                                         
                                                                                                                                     
        global_tmr_voter(1)(548)  <=    (tmr_registers(0)(548) and tmr_registers(1)(548)) or                                            
                            (tmr_registers(1)(548) and tmr_registers(2)(548)) or                                                       
                            (tmr_registers(0)(548) and tmr_registers(2)(548));                                                         
                                                                                                                                     
        global_tmr_voter(1)(549)  <=    (tmr_registers(0)(549) and tmr_registers(1)(549)) or                                            
                            (tmr_registers(1)(549) and tmr_registers(2)(549)) or                                                       
                            (tmr_registers(0)(549) and tmr_registers(2)(549));                                                         
                                                                                                                                     
        global_tmr_voter(1)(550)  <=    (tmr_registers(0)(550) and tmr_registers(1)(550)) or                                            
                            (tmr_registers(1)(550) and tmr_registers(2)(550)) or                                                       
                            (tmr_registers(0)(550) and tmr_registers(2)(550));                                                         
                                                                                                                                     
        global_tmr_voter(1)(551)  <=    (tmr_registers(0)(551) and tmr_registers(1)(551)) or                                            
                            (tmr_registers(1)(551) and tmr_registers(2)(551)) or                                                       
                            (tmr_registers(0)(551) and tmr_registers(2)(551));                                                         
                                                                                                                                     
        global_tmr_voter(1)(552)  <=    (tmr_registers(0)(552) and tmr_registers(1)(552)) or                                            
                            (tmr_registers(1)(552) and tmr_registers(2)(552)) or                                                       
                            (tmr_registers(0)(552) and tmr_registers(2)(552));                                                         
                                                                                                                                     
        global_tmr_voter(1)(553)  <=    (tmr_registers(0)(553) and tmr_registers(1)(553)) or                                            
                            (tmr_registers(1)(553) and tmr_registers(2)(553)) or                                                       
                            (tmr_registers(0)(553) and tmr_registers(2)(553));                                                         
                                                                                                                                     
        global_tmr_voter(1)(554)  <=    (tmr_registers(0)(554) and tmr_registers(1)(554)) or                                            
                            (tmr_registers(1)(554) and tmr_registers(2)(554)) or                                                       
                            (tmr_registers(0)(554) and tmr_registers(2)(554));                                                         
                                                                                                                                     
        global_tmr_voter(1)(555)  <=    (tmr_registers(0)(555) and tmr_registers(1)(555)) or                                            
                            (tmr_registers(1)(555) and tmr_registers(2)(555)) or                                                       
                            (tmr_registers(0)(555) and tmr_registers(2)(555));                                                         
                                                                                                                                     
        global_tmr_voter(1)(556)  <=    (tmr_registers(0)(556) and tmr_registers(1)(556)) or                                            
                            (tmr_registers(1)(556) and tmr_registers(2)(556)) or                                                       
                            (tmr_registers(0)(556) and tmr_registers(2)(556));                                                         
                                                                                                                                     
        global_tmr_voter(1)(557)  <=    (tmr_registers(0)(557) and tmr_registers(1)(557)) or                                            
                            (tmr_registers(1)(557) and tmr_registers(2)(557)) or                                                       
                            (tmr_registers(0)(557) and tmr_registers(2)(557));                                                         
                                                                                                                                     
        global_tmr_voter(1)(558)  <=    (tmr_registers(0)(558) and tmr_registers(1)(558)) or                                            
                            (tmr_registers(1)(558) and tmr_registers(2)(558)) or                                                       
                            (tmr_registers(0)(558) and tmr_registers(2)(558));                                                         
                                                                                                                                     
        global_tmr_voter(1)(559)  <=    (tmr_registers(0)(559) and tmr_registers(1)(559)) or                                            
                            (tmr_registers(1)(559) and tmr_registers(2)(559)) or                                                       
                            (tmr_registers(0)(559) and tmr_registers(2)(559));                                                         
                                                                                                                                     
        global_tmr_voter(1)(560)  <=    (tmr_registers(0)(560) and tmr_registers(1)(560)) or                                            
                            (tmr_registers(1)(560) and tmr_registers(2)(560)) or                                                       
                            (tmr_registers(0)(560) and tmr_registers(2)(560));                                                         
                                                                                                                                     
        global_tmr_voter(1)(561)  <=    (tmr_registers(0)(561) and tmr_registers(1)(561)) or                                            
                            (tmr_registers(1)(561) and tmr_registers(2)(561)) or                                                       
                            (tmr_registers(0)(561) and tmr_registers(2)(561));                                                         
                                                                                                                                     
        global_tmr_voter(1)(562)  <=    (tmr_registers(0)(562) and tmr_registers(1)(562)) or                                            
                            (tmr_registers(1)(562) and tmr_registers(2)(562)) or                                                       
                            (tmr_registers(0)(562) and tmr_registers(2)(562));                                                         
                                                                                                                                     
        global_tmr_voter(1)(563)  <=    (tmr_registers(0)(563) and tmr_registers(1)(563)) or                                            
                            (tmr_registers(1)(563) and tmr_registers(2)(563)) or                                                       
                            (tmr_registers(0)(563) and tmr_registers(2)(563));                                                         
                                                                                                                                     
        global_tmr_voter(1)(564)  <=    (tmr_registers(0)(564) and tmr_registers(1)(564)) or                                            
                            (tmr_registers(1)(564) and tmr_registers(2)(564)) or                                                       
                            (tmr_registers(0)(564) and tmr_registers(2)(564));                                                         
                                                                                                                                     
        global_tmr_voter(1)(565)  <=    (tmr_registers(0)(565) and tmr_registers(1)(565)) or                                            
                            (tmr_registers(1)(565) and tmr_registers(2)(565)) or                                                       
                            (tmr_registers(0)(565) and tmr_registers(2)(565));                                                         
                                                                                                                                     
        global_tmr_voter(1)(566)  <=    (tmr_registers(0)(566) and tmr_registers(1)(566)) or                                            
                            (tmr_registers(1)(566) and tmr_registers(2)(566)) or                                                       
                            (tmr_registers(0)(566) and tmr_registers(2)(566));                                                         
                                                                                                                                     
        global_tmr_voter(1)(567)  <=    (tmr_registers(0)(567) and tmr_registers(1)(567)) or                                            
                            (tmr_registers(1)(567) and tmr_registers(2)(567)) or                                                       
                            (tmr_registers(0)(567) and tmr_registers(2)(567));                                                         
                                                                                                                                     
        global_tmr_voter(1)(568)  <=    (tmr_registers(0)(568) and tmr_registers(1)(568)) or                                            
                            (tmr_registers(1)(568) and tmr_registers(2)(568)) or                                                       
                            (tmr_registers(0)(568) and tmr_registers(2)(568));                                                         
                                                                                                                                     
        global_tmr_voter(1)(569)  <=    (tmr_registers(0)(569) and tmr_registers(1)(569)) or                                            
                            (tmr_registers(1)(569) and tmr_registers(2)(569)) or                                                       
                            (tmr_registers(0)(569) and tmr_registers(2)(569));                                                         
                                                                                                                                     
        global_tmr_voter(1)(570)  <=    (tmr_registers(0)(570) and tmr_registers(1)(570)) or                                            
                            (tmr_registers(1)(570) and tmr_registers(2)(570)) or                                                       
                            (tmr_registers(0)(570) and tmr_registers(2)(570));                                                         
                                                                                                                                     
        global_tmr_voter(1)(571)  <=    (tmr_registers(0)(571) and tmr_registers(1)(571)) or                                            
                            (tmr_registers(1)(571) and tmr_registers(2)(571)) or                                                       
                            (tmr_registers(0)(571) and tmr_registers(2)(571));                                                         
                                                                                                                                     
        global_tmr_voter(1)(572)  <=    (tmr_registers(0)(572) and tmr_registers(1)(572)) or                                            
                            (tmr_registers(1)(572) and tmr_registers(2)(572)) or                                                       
                            (tmr_registers(0)(572) and tmr_registers(2)(572));                                                         
                                                                                                                                     
        global_tmr_voter(1)(573)  <=    (tmr_registers(0)(573) and tmr_registers(1)(573)) or                                            
                            (tmr_registers(1)(573) and tmr_registers(2)(573)) or                                                       
                            (tmr_registers(0)(573) and tmr_registers(2)(573));                                                         
                                                                                                                                     
        global_tmr_voter(1)(574)  <=    (tmr_registers(0)(574) and tmr_registers(1)(574)) or                                            
                            (tmr_registers(1)(574) and tmr_registers(2)(574)) or                                                       
                            (tmr_registers(0)(574) and tmr_registers(2)(574));                                                         
                                                                                                                                     
        global_tmr_voter(1)(575)  <=    (tmr_registers(0)(575) and tmr_registers(1)(575)) or                                            
                            (tmr_registers(1)(575) and tmr_registers(2)(575)) or                                                       
                            (tmr_registers(0)(575) and tmr_registers(2)(575));                                                         
                                                                                                                                     
        global_tmr_voter(1)(576)  <=    (tmr_registers(0)(576) and tmr_registers(1)(576)) or                                            
                            (tmr_registers(1)(576) and tmr_registers(2)(576)) or                                                       
                            (tmr_registers(0)(576) and tmr_registers(2)(576));                                                         
                                                                                                                                     
        global_tmr_voter(1)(577)  <=    (tmr_registers(0)(577) and tmr_registers(1)(577)) or                                            
                            (tmr_registers(1)(577) and tmr_registers(2)(577)) or                                                       
                            (tmr_registers(0)(577) and tmr_registers(2)(577));                                                         
                                                                                                                                     
        global_tmr_voter(1)(578)  <=    (tmr_registers(0)(578) and tmr_registers(1)(578)) or                                            
                            (tmr_registers(1)(578) and tmr_registers(2)(578)) or                                                       
                            (tmr_registers(0)(578) and tmr_registers(2)(578));                                                         
                                                                                                                                     
        global_tmr_voter(1)(579)  <=    (tmr_registers(0)(579) and tmr_registers(1)(579)) or                                            
                            (tmr_registers(1)(579) and tmr_registers(2)(579)) or                                                       
                            (tmr_registers(0)(579) and tmr_registers(2)(579));                                                         
                                                                                                                                     
        global_tmr_voter(1)(580)  <=    (tmr_registers(0)(580) and tmr_registers(1)(580)) or                                            
                            (tmr_registers(1)(580) and tmr_registers(2)(580)) or                                                       
                            (tmr_registers(0)(580) and tmr_registers(2)(580));                                                         
                                                                                                                                     
        global_tmr_voter(1)(581)  <=    (tmr_registers(0)(581) and tmr_registers(1)(581)) or                                            
                            (tmr_registers(1)(581) and tmr_registers(2)(581)) or                                                       
                            (tmr_registers(0)(581) and tmr_registers(2)(581));                                                         
                                                                                                                                     
        global_tmr_voter(1)(582)  <=    (tmr_registers(0)(582) and tmr_registers(1)(582)) or                                            
                            (tmr_registers(1)(582) and tmr_registers(2)(582)) or                                                       
                            (tmr_registers(0)(582) and tmr_registers(2)(582));                                                         
                                                                                                                                     
        global_tmr_voter(1)(583)  <=    (tmr_registers(0)(583) and tmr_registers(1)(583)) or                                            
                            (tmr_registers(1)(583) and tmr_registers(2)(583)) or                                                       
                            (tmr_registers(0)(583) and tmr_registers(2)(583));                                                         
                                                                                                                                     
        global_tmr_voter(1)(584)  <=    (tmr_registers(0)(584) and tmr_registers(1)(584)) or                                            
                            (tmr_registers(1)(584) and tmr_registers(2)(584)) or                                                       
                            (tmr_registers(0)(584) and tmr_registers(2)(584));                                                         
                                                                                                                                     
        global_tmr_voter(1)(585)  <=    (tmr_registers(0)(585) and tmr_registers(1)(585)) or                                            
                            (tmr_registers(1)(585) and tmr_registers(2)(585)) or                                                       
                            (tmr_registers(0)(585) and tmr_registers(2)(585));                                                         
                                                                                                                                     
        global_tmr_voter(1)(586)  <=    (tmr_registers(0)(586) and tmr_registers(1)(586)) or                                            
                            (tmr_registers(1)(586) and tmr_registers(2)(586)) or                                                       
                            (tmr_registers(0)(586) and tmr_registers(2)(586));                                                         
                                                                                                                                     
        global_tmr_voter(1)(587)  <=    (tmr_registers(0)(587) and tmr_registers(1)(587)) or                                            
                            (tmr_registers(1)(587) and tmr_registers(2)(587)) or                                                       
                            (tmr_registers(0)(587) and tmr_registers(2)(587));                                                         
                                                                                                                                     
        global_tmr_voter(1)(588)  <=    (tmr_registers(0)(588) and tmr_registers(1)(588)) or                                            
                            (tmr_registers(1)(588) and tmr_registers(2)(588)) or                                                       
                            (tmr_registers(0)(588) and tmr_registers(2)(588));                                                         
                                                                                                                                     
        global_tmr_voter(1)(589)  <=    (tmr_registers(0)(589) and tmr_registers(1)(589)) or                                            
                            (tmr_registers(1)(589) and tmr_registers(2)(589)) or                                                       
                            (tmr_registers(0)(589) and tmr_registers(2)(589));                                                         
                                                                                                                                     
        global_tmr_voter(1)(590)  <=    (tmr_registers(0)(590) and tmr_registers(1)(590)) or                                            
                            (tmr_registers(1)(590) and tmr_registers(2)(590)) or                                                       
                            (tmr_registers(0)(590) and tmr_registers(2)(590));                                                         
                                                                                                                                     
        global_tmr_voter(1)(591)  <=    (tmr_registers(0)(591) and tmr_registers(1)(591)) or                                            
                            (tmr_registers(1)(591) and tmr_registers(2)(591)) or                                                       
                            (tmr_registers(0)(591) and tmr_registers(2)(591));                                                         
                                                                                                                                     
        global_tmr_voter(1)(592)  <=    (tmr_registers(0)(592) and tmr_registers(1)(592)) or                                            
                            (tmr_registers(1)(592) and tmr_registers(2)(592)) or                                                       
                            (tmr_registers(0)(592) and tmr_registers(2)(592));                                                         
                                                                                                                                     
        global_tmr_voter(1)(593)  <=    (tmr_registers(0)(593) and tmr_registers(1)(593)) or                                            
                            (tmr_registers(1)(593) and tmr_registers(2)(593)) or                                                       
                            (tmr_registers(0)(593) and tmr_registers(2)(593));                                                         
                                                                                                                                     
        global_tmr_voter(1)(594)  <=    (tmr_registers(0)(594) and tmr_registers(1)(594)) or                                            
                            (tmr_registers(1)(594) and tmr_registers(2)(594)) or                                                       
                            (tmr_registers(0)(594) and tmr_registers(2)(594));                                                         
                                                                                                                                     
        global_tmr_voter(1)(595)  <=    (tmr_registers(0)(595) and tmr_registers(1)(595)) or                                            
                            (tmr_registers(1)(595) and tmr_registers(2)(595)) or                                                       
                            (tmr_registers(0)(595) and tmr_registers(2)(595));                                                         
                                                                                                                                     
        global_tmr_voter(1)(596)  <=    (tmr_registers(0)(596) and tmr_registers(1)(596)) or                                            
                            (tmr_registers(1)(596) and tmr_registers(2)(596)) or                                                       
                            (tmr_registers(0)(596) and tmr_registers(2)(596));                                                         
                                                                                                                                     
        global_tmr_voter(1)(597)  <=    (tmr_registers(0)(597) and tmr_registers(1)(597)) or                                            
                            (tmr_registers(1)(597) and tmr_registers(2)(597)) or                                                       
                            (tmr_registers(0)(597) and tmr_registers(2)(597));                                                         
                                                                                                                                     
        global_tmr_voter(1)(598)  <=    (tmr_registers(0)(598) and tmr_registers(1)(598)) or                                            
                            (tmr_registers(1)(598) and tmr_registers(2)(598)) or                                                       
                            (tmr_registers(0)(598) and tmr_registers(2)(598));                                                         
                                                                                                                                     
        global_tmr_voter(1)(599)  <=    (tmr_registers(0)(599) and tmr_registers(1)(599)) or                                            
                            (tmr_registers(1)(599) and tmr_registers(2)(599)) or                                                       
                            (tmr_registers(0)(599) and tmr_registers(2)(599));                                                         
                                                                                                                                     
        global_tmr_voter(1)(600)  <=    (tmr_registers(0)(600) and tmr_registers(1)(600)) or                                            
                            (tmr_registers(1)(600) and tmr_registers(2)(600)) or                                                       
                            (tmr_registers(0)(600) and tmr_registers(2)(600));                                                         
                                                                                                                                     
        global_tmr_voter(1)(601)  <=    (tmr_registers(0)(601) and tmr_registers(1)(601)) or                                            
                            (tmr_registers(1)(601) and tmr_registers(2)(601)) or                                                       
                            (tmr_registers(0)(601) and tmr_registers(2)(601));                                                         
                                                                                                                                     
        global_tmr_voter(1)(602)  <=    (tmr_registers(0)(602) and tmr_registers(1)(602)) or                                            
                            (tmr_registers(1)(602) and tmr_registers(2)(602)) or                                                       
                            (tmr_registers(0)(602) and tmr_registers(2)(602));                                                         
                                                                                                                                     
        global_tmr_voter(1)(603)  <=    (tmr_registers(0)(603) and tmr_registers(1)(603)) or                                            
                            (tmr_registers(1)(603) and tmr_registers(2)(603)) or                                                       
                            (tmr_registers(0)(603) and tmr_registers(2)(603));                                                         
                                                                                                                                     
        global_tmr_voter(1)(604)  <=    (tmr_registers(0)(604) and tmr_registers(1)(604)) or                                            
                            (tmr_registers(1)(604) and tmr_registers(2)(604)) or                                                       
                            (tmr_registers(0)(604) and tmr_registers(2)(604));                                                         
                                                                                                                                     
        global_tmr_voter(1)(605)  <=    (tmr_registers(0)(605) and tmr_registers(1)(605)) or                                            
                            (tmr_registers(1)(605) and tmr_registers(2)(605)) or                                                       
                            (tmr_registers(0)(605) and tmr_registers(2)(605));                                                         
                                                                                                                                     
        global_tmr_voter(1)(606)  <=    (tmr_registers(0)(606) and tmr_registers(1)(606)) or                                            
                            (tmr_registers(1)(606) and tmr_registers(2)(606)) or                                                       
                            (tmr_registers(0)(606) and tmr_registers(2)(606));                                                         
                                                                                                                                     
        global_tmr_voter(1)(607)  <=    (tmr_registers(0)(607) and tmr_registers(1)(607)) or                                            
                            (tmr_registers(1)(607) and tmr_registers(2)(607)) or                                                       
                            (tmr_registers(0)(607) and tmr_registers(2)(607));                                                         
                                                                                                                                     
        global_tmr_voter(1)(608)  <=    (tmr_registers(0)(608) and tmr_registers(1)(608)) or                                            
                            (tmr_registers(1)(608) and tmr_registers(2)(608)) or                                                       
                            (tmr_registers(0)(608) and tmr_registers(2)(608));                                                         
                                                                                                                                     
        global_tmr_voter(1)(609)  <=    (tmr_registers(0)(609) and tmr_registers(1)(609)) or                                            
                            (tmr_registers(1)(609) and tmr_registers(2)(609)) or                                                       
                            (tmr_registers(0)(609) and tmr_registers(2)(609));                                                         
                                                                                                                                     
        global_tmr_voter(1)(610)  <=    (tmr_registers(0)(610) and tmr_registers(1)(610)) or                                            
                            (tmr_registers(1)(610) and tmr_registers(2)(610)) or                                                       
                            (tmr_registers(0)(610) and tmr_registers(2)(610));                                                         
                                                                                                                                     
        global_tmr_voter(1)(611)  <=    (tmr_registers(0)(611) and tmr_registers(1)(611)) or                                            
                            (tmr_registers(1)(611) and tmr_registers(2)(611)) or                                                       
                            (tmr_registers(0)(611) and tmr_registers(2)(611));                                                         
                                                                                                                                     
        global_tmr_voter(1)(612)  <=    (tmr_registers(0)(612) and tmr_registers(1)(612)) or                                            
                            (tmr_registers(1)(612) and tmr_registers(2)(612)) or                                                       
                            (tmr_registers(0)(612) and tmr_registers(2)(612));                                                         
                                                                                                                                     
        global_tmr_voter(1)(613)  <=    (tmr_registers(0)(613) and tmr_registers(1)(613)) or                                            
                            (tmr_registers(1)(613) and tmr_registers(2)(613)) or                                                       
                            (tmr_registers(0)(613) and tmr_registers(2)(613));                                                         
                                                                                                                                     
        global_tmr_voter(1)(614)  <=    (tmr_registers(0)(614) and tmr_registers(1)(614)) or                                            
                            (tmr_registers(1)(614) and tmr_registers(2)(614)) or                                                       
                            (tmr_registers(0)(614) and tmr_registers(2)(614));                                                         
                                                                                                                                     
        global_tmr_voter(1)(615)  <=    (tmr_registers(0)(615) and tmr_registers(1)(615)) or                                            
                            (tmr_registers(1)(615) and tmr_registers(2)(615)) or                                                       
                            (tmr_registers(0)(615) and tmr_registers(2)(615));                                                         
                                                                                                                                     
        global_tmr_voter(1)(616)  <=    (tmr_registers(0)(616) and tmr_registers(1)(616)) or                                            
                            (tmr_registers(1)(616) and tmr_registers(2)(616)) or                                                       
                            (tmr_registers(0)(616) and tmr_registers(2)(616));                                                         
                                                                                                                                     
        global_tmr_voter(1)(617)  <=    (tmr_registers(0)(617) and tmr_registers(1)(617)) or                                            
                            (tmr_registers(1)(617) and tmr_registers(2)(617)) or                                                       
                            (tmr_registers(0)(617) and tmr_registers(2)(617));                                                         
                                                                                                                                     
        global_tmr_voter(1)(618)  <=    (tmr_registers(0)(618) and tmr_registers(1)(618)) or                                            
                            (tmr_registers(1)(618) and tmr_registers(2)(618)) or                                                       
                            (tmr_registers(0)(618) and tmr_registers(2)(618));                                                         
                                                                                                                                     
        global_tmr_voter(1)(619)  <=    (tmr_registers(0)(619) and tmr_registers(1)(619)) or                                            
                            (tmr_registers(1)(619) and tmr_registers(2)(619)) or                                                       
                            (tmr_registers(0)(619) and tmr_registers(2)(619));                                                         
                                                                                                                                     
        global_tmr_voter(1)(620)  <=    (tmr_registers(0)(620) and tmr_registers(1)(620)) or                                            
                            (tmr_registers(1)(620) and tmr_registers(2)(620)) or                                                       
                            (tmr_registers(0)(620) and tmr_registers(2)(620));                                                         
                                                                                                                                     
        global_tmr_voter(1)(621)  <=    (tmr_registers(0)(621) and tmr_registers(1)(621)) or                                            
                            (tmr_registers(1)(621) and tmr_registers(2)(621)) or                                                       
                            (tmr_registers(0)(621) and tmr_registers(2)(621));                                                         
                                                                                                                                     
        global_tmr_voter(1)(622)  <=    (tmr_registers(0)(622) and tmr_registers(1)(622)) or                                            
                            (tmr_registers(1)(622) and tmr_registers(2)(622)) or                                                       
                            (tmr_registers(0)(622) and tmr_registers(2)(622));                                                         
                                                                                                                                     
        global_tmr_voter(1)(623)  <=    (tmr_registers(0)(623) and tmr_registers(1)(623)) or                                            
                            (tmr_registers(1)(623) and tmr_registers(2)(623)) or                                                       
                            (tmr_registers(0)(623) and tmr_registers(2)(623));                                                         
                                                                                                                                     
        global_tmr_voter(1)(624)  <=    (tmr_registers(0)(624) and tmr_registers(1)(624)) or                                            
                            (tmr_registers(1)(624) and tmr_registers(2)(624)) or                                                       
                            (tmr_registers(0)(624) and tmr_registers(2)(624));                                                         
                                                                                                                                     
        global_tmr_voter(1)(625)  <=    (tmr_registers(0)(625) and tmr_registers(1)(625)) or                                            
                            (tmr_registers(1)(625) and tmr_registers(2)(625)) or                                                       
                            (tmr_registers(0)(625) and tmr_registers(2)(625));                                                         
                                                                                                                                     
        global_tmr_voter(1)(626)  <=    (tmr_registers(0)(626) and tmr_registers(1)(626)) or                                            
                            (tmr_registers(1)(626) and tmr_registers(2)(626)) or                                                       
                            (tmr_registers(0)(626) and tmr_registers(2)(626));                                                         
                                                                                                                                     
        global_tmr_voter(1)(627)  <=    (tmr_registers(0)(627) and tmr_registers(1)(627)) or                                            
                            (tmr_registers(1)(627) and tmr_registers(2)(627)) or                                                       
                            (tmr_registers(0)(627) and tmr_registers(2)(627));                                                         
                                                                                                                                     
        global_tmr_voter(1)(628)  <=    (tmr_registers(0)(628) and tmr_registers(1)(628)) or                                            
                            (tmr_registers(1)(628) and tmr_registers(2)(628)) or                                                       
                            (tmr_registers(0)(628) and tmr_registers(2)(628));                                                         
                                                                                                                                     
        global_tmr_voter(1)(629)  <=    (tmr_registers(0)(629) and tmr_registers(1)(629)) or                                            
                            (tmr_registers(1)(629) and tmr_registers(2)(629)) or                                                       
                            (tmr_registers(0)(629) and tmr_registers(2)(629));                                                         
                                                                                                                                     
        global_tmr_voter(1)(630)  <=    (tmr_registers(0)(630) and tmr_registers(1)(630)) or                                            
                            (tmr_registers(1)(630) and tmr_registers(2)(630)) or                                                       
                            (tmr_registers(0)(630) and tmr_registers(2)(630));                                                         
                                                                                                                                     
        global_tmr_voter(1)(631)  <=    (tmr_registers(0)(631) and tmr_registers(1)(631)) or                                            
                            (tmr_registers(1)(631) and tmr_registers(2)(631)) or                                                       
                            (tmr_registers(0)(631) and tmr_registers(2)(631));                                                         
                                                                                                                                     
        global_tmr_voter(1)(632)  <=    (tmr_registers(0)(632) and tmr_registers(1)(632)) or                                            
                            (tmr_registers(1)(632) and tmr_registers(2)(632)) or                                                       
                            (tmr_registers(0)(632) and tmr_registers(2)(632));                                                         
                                                                                                                                     
        global_tmr_voter(1)(633)  <=    (tmr_registers(0)(633) and tmr_registers(1)(633)) or                                            
                            (tmr_registers(1)(633) and tmr_registers(2)(633)) or                                                       
                            (tmr_registers(0)(633) and tmr_registers(2)(633));                                                         
                                                                                                                                     
        global_tmr_voter(1)(634)  <=    (tmr_registers(0)(634) and tmr_registers(1)(634)) or                                            
                            (tmr_registers(1)(634) and tmr_registers(2)(634)) or                                                       
                            (tmr_registers(0)(634) and tmr_registers(2)(634));                                                         
                                                                                                                                     
        global_tmr_voter(1)(635)  <=    (tmr_registers(0)(635) and tmr_registers(1)(635)) or                                            
                            (tmr_registers(1)(635) and tmr_registers(2)(635)) or                                                       
                            (tmr_registers(0)(635) and tmr_registers(2)(635));                                                         
                                                                                                                                     
        global_tmr_voter(1)(636)  <=    (tmr_registers(0)(636) and tmr_registers(1)(636)) or                                            
                            (tmr_registers(1)(636) and tmr_registers(2)(636)) or                                                       
                            (tmr_registers(0)(636) and tmr_registers(2)(636));                                                         
                                                                                                                                     
        global_tmr_voter(1)(637)  <=    (tmr_registers(0)(637) and tmr_registers(1)(637)) or                                            
                            (tmr_registers(1)(637) and tmr_registers(2)(637)) or                                                       
                            (tmr_registers(0)(637) and tmr_registers(2)(637));                                                         
                                                                                                                                     
        global_tmr_voter(1)(638)  <=    (tmr_registers(0)(638) and tmr_registers(1)(638)) or                                            
                            (tmr_registers(1)(638) and tmr_registers(2)(638)) or                                                       
                            (tmr_registers(0)(638) and tmr_registers(2)(638));                                                         
                                                                                                                                     
        global_tmr_voter(1)(639)  <=    (tmr_registers(0)(639) and tmr_registers(1)(639)) or                                            
                            (tmr_registers(1)(639) and tmr_registers(2)(639)) or                                                       
                            (tmr_registers(0)(639) and tmr_registers(2)(639));                                                         
                                                                                                                                     
        global_tmr_voter(1)(640)  <=    (tmr_registers(0)(640) and tmr_registers(1)(640)) or                                            
                            (tmr_registers(1)(640) and tmr_registers(2)(640)) or                                                       
                            (tmr_registers(0)(640) and tmr_registers(2)(640));                                                         
                                                                                                                                     
        global_tmr_voter(1)(641)  <=    (tmr_registers(0)(641) and tmr_registers(1)(641)) or                                            
                            (tmr_registers(1)(641) and tmr_registers(2)(641)) or                                                       
                            (tmr_registers(0)(641) and tmr_registers(2)(641));                                                         
                                                                                                                                     
        global_tmr_voter(1)(642)  <=    (tmr_registers(0)(642) and tmr_registers(1)(642)) or                                            
                            (tmr_registers(1)(642) and tmr_registers(2)(642)) or                                                       
                            (tmr_registers(0)(642) and tmr_registers(2)(642));                                                         
                                                                                                                                     
        global_tmr_voter(1)(643)  <=    (tmr_registers(0)(643) and tmr_registers(1)(643)) or                                            
                            (tmr_registers(1)(643) and tmr_registers(2)(643)) or                                                       
                            (tmr_registers(0)(643) and tmr_registers(2)(643));                                                         
                                                                                                                                     
        global_tmr_voter(1)(644)  <=    (tmr_registers(0)(644) and tmr_registers(1)(644)) or                                            
                            (tmr_registers(1)(644) and tmr_registers(2)(644)) or                                                       
                            (tmr_registers(0)(644) and tmr_registers(2)(644));                                                         
                                                                                                                                     
        global_tmr_voter(1)(645)  <=    (tmr_registers(0)(645) and tmr_registers(1)(645)) or                                            
                            (tmr_registers(1)(645) and tmr_registers(2)(645)) or                                                       
                            (tmr_registers(0)(645) and tmr_registers(2)(645));                                                         
                                                                                                                                     
        global_tmr_voter(1)(646)  <=    (tmr_registers(0)(646) and tmr_registers(1)(646)) or                                            
                            (tmr_registers(1)(646) and tmr_registers(2)(646)) or                                                       
                            (tmr_registers(0)(646) and tmr_registers(2)(646));                                                         
                                                                                                                                     
        global_tmr_voter(1)(647)  <=    (tmr_registers(0)(647) and tmr_registers(1)(647)) or                                            
                            (tmr_registers(1)(647) and tmr_registers(2)(647)) or                                                       
                            (tmr_registers(0)(647) and tmr_registers(2)(647));                                                         
                                                                                                                                     
        global_tmr_voter(1)(648)  <=    (tmr_registers(0)(648) and tmr_registers(1)(648)) or                                            
                            (tmr_registers(1)(648) and tmr_registers(2)(648)) or                                                       
                            (tmr_registers(0)(648) and tmr_registers(2)(648));                                                         
                                                                                                                                     
        global_tmr_voter(1)(649)  <=    (tmr_registers(0)(649) and tmr_registers(1)(649)) or                                            
                            (tmr_registers(1)(649) and tmr_registers(2)(649)) or                                                       
                            (tmr_registers(0)(649) and tmr_registers(2)(649));                                                         
                                                                                                                                     
        global_tmr_voter(1)(650)  <=    (tmr_registers(0)(650) and tmr_registers(1)(650)) or                                            
                            (tmr_registers(1)(650) and tmr_registers(2)(650)) or                                                       
                            (tmr_registers(0)(650) and tmr_registers(2)(650));                                                         
                                                                                                                                     
        global_tmr_voter(1)(651)  <=    (tmr_registers(0)(651) and tmr_registers(1)(651)) or                                            
                            (tmr_registers(1)(651) and tmr_registers(2)(651)) or                                                       
                            (tmr_registers(0)(651) and tmr_registers(2)(651));                                                         
                                                                                                                                     
        global_tmr_voter(1)(652)  <=    (tmr_registers(0)(652) and tmr_registers(1)(652)) or                                            
                            (tmr_registers(1)(652) and tmr_registers(2)(652)) or                                                       
                            (tmr_registers(0)(652) and tmr_registers(2)(652));                                                         
                                                                                                                                     
        global_tmr_voter(1)(653)  <=    (tmr_registers(0)(653) and tmr_registers(1)(653)) or                                            
                            (tmr_registers(1)(653) and tmr_registers(2)(653)) or                                                       
                            (tmr_registers(0)(653) and tmr_registers(2)(653));                                                         
                                                                                                                                     
        global_tmr_voter(1)(654)  <=    (tmr_registers(0)(654) and tmr_registers(1)(654)) or                                            
                            (tmr_registers(1)(654) and tmr_registers(2)(654)) or                                                       
                            (tmr_registers(0)(654) and tmr_registers(2)(654));                                                         
                                                                                                                                     
        global_tmr_voter(1)(655)  <=    (tmr_registers(0)(655) and tmr_registers(1)(655)) or                                            
                            (tmr_registers(1)(655) and tmr_registers(2)(655)) or                                                       
                            (tmr_registers(0)(655) and tmr_registers(2)(655));                                                         
                                                                                                                                     
        global_tmr_voter(1)(656)  <=    (tmr_registers(0)(656) and tmr_registers(1)(656)) or                                            
                            (tmr_registers(1)(656) and tmr_registers(2)(656)) or                                                       
                            (tmr_registers(0)(656) and tmr_registers(2)(656));                                                         
                                                                                                                                     
        global_tmr_voter(1)(657)  <=    (tmr_registers(0)(657) and tmr_registers(1)(657)) or                                            
                            (tmr_registers(1)(657) and tmr_registers(2)(657)) or                                                       
                            (tmr_registers(0)(657) and tmr_registers(2)(657));                                                         
                                                                                                                                     
        global_tmr_voter(1)(658)  <=    (tmr_registers(0)(658) and tmr_registers(1)(658)) or                                            
                            (tmr_registers(1)(658) and tmr_registers(2)(658)) or                                                       
                            (tmr_registers(0)(658) and tmr_registers(2)(658));                                                         
                                                                                                                                     
        global_tmr_voter(1)(659)  <=    (tmr_registers(0)(659) and tmr_registers(1)(659)) or                                            
                            (tmr_registers(1)(659) and tmr_registers(2)(659)) or                                                       
                            (tmr_registers(0)(659) and tmr_registers(2)(659));                                                         
                                                                                                                                     
        global_tmr_voter(1)(660)  <=    (tmr_registers(0)(660) and tmr_registers(1)(660)) or                                            
                            (tmr_registers(1)(660) and tmr_registers(2)(660)) or                                                       
                            (tmr_registers(0)(660) and tmr_registers(2)(660));                                                         
                                                                                                                                     
        global_tmr_voter(1)(661)  <=    (tmr_registers(0)(661) and tmr_registers(1)(661)) or                                            
                            (tmr_registers(1)(661) and tmr_registers(2)(661)) or                                                       
                            (tmr_registers(0)(661) and tmr_registers(2)(661));                                                         
                                                                                                                                     
        global_tmr_voter(1)(662)  <=    (tmr_registers(0)(662) and tmr_registers(1)(662)) or                                            
                            (tmr_registers(1)(662) and tmr_registers(2)(662)) or                                                       
                            (tmr_registers(0)(662) and tmr_registers(2)(662));                                                         
                                                                                                                                     
        global_tmr_voter(1)(663)  <=    (tmr_registers(0)(663) and tmr_registers(1)(663)) or                                            
                            (tmr_registers(1)(663) and tmr_registers(2)(663)) or                                                       
                            (tmr_registers(0)(663) and tmr_registers(2)(663));                                                         
                                                                                                                                     
        global_tmr_voter(1)(664)  <=    (tmr_registers(0)(664) and tmr_registers(1)(664)) or                                            
                            (tmr_registers(1)(664) and tmr_registers(2)(664)) or                                                       
                            (tmr_registers(0)(664) and tmr_registers(2)(664));                                                         
                                                                                                                                     
        global_tmr_voter(1)(665)  <=    (tmr_registers(0)(665) and tmr_registers(1)(665)) or                                            
                            (tmr_registers(1)(665) and tmr_registers(2)(665)) or                                                       
                            (tmr_registers(0)(665) and tmr_registers(2)(665));                                                         
                                                                                                                                     
        global_tmr_voter(1)(666)  <=    (tmr_registers(0)(666) and tmr_registers(1)(666)) or                                            
                            (tmr_registers(1)(666) and tmr_registers(2)(666)) or                                                       
                            (tmr_registers(0)(666) and tmr_registers(2)(666));                                                         
                                                                                                                                     
        global_tmr_voter(1)(667)  <=    (tmr_registers(0)(667) and tmr_registers(1)(667)) or                                            
                            (tmr_registers(1)(667) and tmr_registers(2)(667)) or                                                       
                            (tmr_registers(0)(667) and tmr_registers(2)(667));                                                         
                                                                                                                                     
        global_tmr_voter(1)(668)  <=    (tmr_registers(0)(668) and tmr_registers(1)(668)) or                                            
                            (tmr_registers(1)(668) and tmr_registers(2)(668)) or                                                       
                            (tmr_registers(0)(668) and tmr_registers(2)(668));                                                         
                                                                                                                                     
        global_tmr_voter(1)(669)  <=    (tmr_registers(0)(669) and tmr_registers(1)(669)) or                                            
                            (tmr_registers(1)(669) and tmr_registers(2)(669)) or                                                       
                            (tmr_registers(0)(669) and tmr_registers(2)(669));                                                         
                                                                                                                                     
        global_tmr_voter(1)(670)  <=    (tmr_registers(0)(670) and tmr_registers(1)(670)) or                                            
                            (tmr_registers(1)(670) and tmr_registers(2)(670)) or                                                       
                            (tmr_registers(0)(670) and tmr_registers(2)(670));                                                         
                                                                                                                                     
        global_tmr_voter(1)(671)  <=    (tmr_registers(0)(671) and tmr_registers(1)(671)) or                                            
                            (tmr_registers(1)(671) and tmr_registers(2)(671)) or                                                       
                            (tmr_registers(0)(671) and tmr_registers(2)(671));                                                         
                                                                                                                                     
        global_tmr_voter(1)(672)  <=    (tmr_registers(0)(672) and tmr_registers(1)(672)) or                                            
                            (tmr_registers(1)(672) and tmr_registers(2)(672)) or                                                       
                            (tmr_registers(0)(672) and tmr_registers(2)(672));                                                         
                                                                                                                                     
        global_tmr_voter(1)(673)  <=    (tmr_registers(0)(673) and tmr_registers(1)(673)) or                                            
                            (tmr_registers(1)(673) and tmr_registers(2)(673)) or                                                       
                            (tmr_registers(0)(673) and tmr_registers(2)(673));                                                         
                                                                                                                                     
        global_tmr_voter(1)(674)  <=    (tmr_registers(0)(674) and tmr_registers(1)(674)) or                                            
                            (tmr_registers(1)(674) and tmr_registers(2)(674)) or                                                       
                            (tmr_registers(0)(674) and tmr_registers(2)(674));                                                         
                                                                                                                                     
        global_tmr_voter(1)(675)  <=    (tmr_registers(0)(675) and tmr_registers(1)(675)) or                                            
                            (tmr_registers(1)(675) and tmr_registers(2)(675)) or                                                       
                            (tmr_registers(0)(675) and tmr_registers(2)(675));                                                         
                                                                                                                                     
        global_tmr_voter(1)(676)  <=    (tmr_registers(0)(676) and tmr_registers(1)(676)) or                                            
                            (tmr_registers(1)(676) and tmr_registers(2)(676)) or                                                       
                            (tmr_registers(0)(676) and tmr_registers(2)(676));                                                         
                                                                                                                                     
        global_tmr_voter(1)(677)  <=    (tmr_registers(0)(677) and tmr_registers(1)(677)) or                                            
                            (tmr_registers(1)(677) and tmr_registers(2)(677)) or                                                       
                            (tmr_registers(0)(677) and tmr_registers(2)(677));                                                         
                                                                                                                                     
        global_tmr_voter(1)(678)  <=    (tmr_registers(0)(678) and tmr_registers(1)(678)) or                                            
                            (tmr_registers(1)(678) and tmr_registers(2)(678)) or                                                       
                            (tmr_registers(0)(678) and tmr_registers(2)(678));                                                         
                                                                                                                                     
        global_tmr_voter(1)(679)  <=    (tmr_registers(0)(679) and tmr_registers(1)(679)) or                                            
                            (tmr_registers(1)(679) and tmr_registers(2)(679)) or                                                       
                            (tmr_registers(0)(679) and tmr_registers(2)(679));                                                         
                                                                                                                                     
        global_tmr_voter(1)(680)  <=    (tmr_registers(0)(680) and tmr_registers(1)(680)) or                                            
                            (tmr_registers(1)(680) and tmr_registers(2)(680)) or                                                       
                            (tmr_registers(0)(680) and tmr_registers(2)(680));                                                         
                                                                                                                                     
        global_tmr_voter(1)(681)  <=    (tmr_registers(0)(681) and tmr_registers(1)(681)) or                                            
                            (tmr_registers(1)(681) and tmr_registers(2)(681)) or                                                       
                            (tmr_registers(0)(681) and tmr_registers(2)(681));                                                         
                                                                                                                                     
        global_tmr_voter(1)(682)  <=    (tmr_registers(0)(682) and tmr_registers(1)(682)) or                                            
                            (tmr_registers(1)(682) and tmr_registers(2)(682)) or                                                       
                            (tmr_registers(0)(682) and tmr_registers(2)(682));                                                         
                                                                                                                                     
        global_tmr_voter(1)(683)  <=    (tmr_registers(0)(683) and tmr_registers(1)(683)) or                                            
                            (tmr_registers(1)(683) and tmr_registers(2)(683)) or                                                       
                            (tmr_registers(0)(683) and tmr_registers(2)(683));                                                         
                                                                                                                                     
        global_tmr_voter(1)(684)  <=    (tmr_registers(0)(684) and tmr_registers(1)(684)) or                                            
                            (tmr_registers(1)(684) and tmr_registers(2)(684)) or                                                       
                            (tmr_registers(0)(684) and tmr_registers(2)(684));                                                         
                                                                                                                                     
        global_tmr_voter(1)(685)  <=    (tmr_registers(0)(685) and tmr_registers(1)(685)) or                                            
                            (tmr_registers(1)(685) and tmr_registers(2)(685)) or                                                       
                            (tmr_registers(0)(685) and tmr_registers(2)(685));                                                         
                                                                                                                                     
        global_tmr_voter(1)(686)  <=    (tmr_registers(0)(686) and tmr_registers(1)(686)) or                                            
                            (tmr_registers(1)(686) and tmr_registers(2)(686)) or                                                       
                            (tmr_registers(0)(686) and tmr_registers(2)(686));                                                         
                                                                                                                                     
        global_tmr_voter(1)(687)  <=    (tmr_registers(0)(687) and tmr_registers(1)(687)) or                                            
                            (tmr_registers(1)(687) and tmr_registers(2)(687)) or                                                       
                            (tmr_registers(0)(687) and tmr_registers(2)(687));                                                         
                                                                                                                                     
        global_tmr_voter(1)(688)  <=    (tmr_registers(0)(688) and tmr_registers(1)(688)) or                                            
                            (tmr_registers(1)(688) and tmr_registers(2)(688)) or                                                       
                            (tmr_registers(0)(688) and tmr_registers(2)(688));                                                         
                                                                                                                                     
        global_tmr_voter(1)(689)  <=    (tmr_registers(0)(689) and tmr_registers(1)(689)) or                                            
                            (tmr_registers(1)(689) and tmr_registers(2)(689)) or                                                       
                            (tmr_registers(0)(689) and tmr_registers(2)(689));                                                         
                                                                                                                                     
        global_tmr_voter(1)(690)  <=    (tmr_registers(0)(690) and tmr_registers(1)(690)) or                                            
                            (tmr_registers(1)(690) and tmr_registers(2)(690)) or                                                       
                            (tmr_registers(0)(690) and tmr_registers(2)(690));                                                         
                                                                                                                                     
        global_tmr_voter(1)(691)  <=    (tmr_registers(0)(691) and tmr_registers(1)(691)) or                                            
                            (tmr_registers(1)(691) and tmr_registers(2)(691)) or                                                       
                            (tmr_registers(0)(691) and tmr_registers(2)(691));                                                         
                                                                                                                                     
        global_tmr_voter(1)(692)  <=    (tmr_registers(0)(692) and tmr_registers(1)(692)) or                                            
                            (tmr_registers(1)(692) and tmr_registers(2)(692)) or                                                       
                            (tmr_registers(0)(692) and tmr_registers(2)(692));                                                         
                                                                                                                                     
        global_tmr_voter(1)(693)  <=    (tmr_registers(0)(693) and tmr_registers(1)(693)) or                                            
                            (tmr_registers(1)(693) and tmr_registers(2)(693)) or                                                       
                            (tmr_registers(0)(693) and tmr_registers(2)(693));                                                         
                                                                                                                                     
        global_tmr_voter(1)(694)  <=    (tmr_registers(0)(694) and tmr_registers(1)(694)) or                                            
                            (tmr_registers(1)(694) and tmr_registers(2)(694)) or                                                       
                            (tmr_registers(0)(694) and tmr_registers(2)(694));                                                         
                                                                                                                                     
        global_tmr_voter(1)(695)  <=    (tmr_registers(0)(695) and tmr_registers(1)(695)) or                                            
                            (tmr_registers(1)(695) and tmr_registers(2)(695)) or                                                       
                            (tmr_registers(0)(695) and tmr_registers(2)(695));                                                         
                                                                                                                                     
        global_tmr_voter(1)(696)  <=    (tmr_registers(0)(696) and tmr_registers(1)(696)) or                                            
                            (tmr_registers(1)(696) and tmr_registers(2)(696)) or                                                       
                            (tmr_registers(0)(696) and tmr_registers(2)(696));                                                         
                                                                                                                                     
        global_tmr_voter(1)(697)  <=    (tmr_registers(0)(697) and tmr_registers(1)(697)) or                                            
                            (tmr_registers(1)(697) and tmr_registers(2)(697)) or                                                       
                            (tmr_registers(0)(697) and tmr_registers(2)(697));                                                         
                                                                                                                                     
        global_tmr_voter(1)(698)  <=    (tmr_registers(0)(698) and tmr_registers(1)(698)) or                                            
                            (tmr_registers(1)(698) and tmr_registers(2)(698)) or                                                       
                            (tmr_registers(0)(698) and tmr_registers(2)(698));                                                         
                                                                                                                                     
        global_tmr_voter(1)(699)  <=    (tmr_registers(0)(699) and tmr_registers(1)(699)) or                                            
                            (tmr_registers(1)(699) and tmr_registers(2)(699)) or                                                       
                            (tmr_registers(0)(699) and tmr_registers(2)(699));                                                         
                                                                                                                                     
        global_tmr_voter(1)(700)  <=    (tmr_registers(0)(700) and tmr_registers(1)(700)) or                                            
                            (tmr_registers(1)(700) and tmr_registers(2)(700)) or                                                       
                            (tmr_registers(0)(700) and tmr_registers(2)(700));                                                         
                                                                                                                                     
        global_tmr_voter(1)(701)  <=    (tmr_registers(0)(701) and tmr_registers(1)(701)) or                                            
                            (tmr_registers(1)(701) and tmr_registers(2)(701)) or                                                       
                            (tmr_registers(0)(701) and tmr_registers(2)(701));                                                         
                                                                                                                                     
        global_tmr_voter(1)(702)  <=    (tmr_registers(0)(702) and tmr_registers(1)(702)) or                                            
                            (tmr_registers(1)(702) and tmr_registers(2)(702)) or                                                       
                            (tmr_registers(0)(702) and tmr_registers(2)(702));                                                         
                                                                                                                                     
        global_tmr_voter(1)(703)  <=    (tmr_registers(0)(703) and tmr_registers(1)(703)) or                                            
                            (tmr_registers(1)(703) and tmr_registers(2)(703)) or                                                       
                            (tmr_registers(0)(703) and tmr_registers(2)(703));                                                         
                                                                                                                                     
        global_tmr_voter(1)(704)  <=    (tmr_registers(0)(704) and tmr_registers(1)(704)) or                                            
                            (tmr_registers(1)(704) and tmr_registers(2)(704)) or                                                       
                            (tmr_registers(0)(704) and tmr_registers(2)(704));                                                         
                                                                                                                                     
        global_tmr_voter(1)(705)  <=    (tmr_registers(0)(705) and tmr_registers(1)(705)) or                                            
                            (tmr_registers(1)(705) and tmr_registers(2)(705)) or                                                       
                            (tmr_registers(0)(705) and tmr_registers(2)(705));                                                         
                                                                                                                                     
        global_tmr_voter(1)(706)  <=    (tmr_registers(0)(706) and tmr_registers(1)(706)) or                                            
                            (tmr_registers(1)(706) and tmr_registers(2)(706)) or                                                       
                            (tmr_registers(0)(706) and tmr_registers(2)(706));                                                         
                                                                                                                                     
        global_tmr_voter(1)(707)  <=    (tmr_registers(0)(707) and tmr_registers(1)(707)) or                                            
                            (tmr_registers(1)(707) and tmr_registers(2)(707)) or                                                       
                            (tmr_registers(0)(707) and tmr_registers(2)(707));                                                         
                                                                                                                                     
        global_tmr_voter(1)(708)  <=    (tmr_registers(0)(708) and tmr_registers(1)(708)) or                                            
                            (tmr_registers(1)(708) and tmr_registers(2)(708)) or                                                       
                            (tmr_registers(0)(708) and tmr_registers(2)(708));                                                         
                                                                                                                                     
        global_tmr_voter(1)(709)  <=    (tmr_registers(0)(709) and tmr_registers(1)(709)) or                                            
                            (tmr_registers(1)(709) and tmr_registers(2)(709)) or                                                       
                            (tmr_registers(0)(709) and tmr_registers(2)(709));                                                         
                                                                                                                                     
        global_tmr_voter(1)(710)  <=    (tmr_registers(0)(710) and tmr_registers(1)(710)) or                                            
                            (tmr_registers(1)(710) and tmr_registers(2)(710)) or                                                       
                            (tmr_registers(0)(710) and tmr_registers(2)(710));                                                         
                                                                                                                                     
        global_tmr_voter(1)(711)  <=    (tmr_registers(0)(711) and tmr_registers(1)(711)) or                                            
                            (tmr_registers(1)(711) and tmr_registers(2)(711)) or                                                       
                            (tmr_registers(0)(711) and tmr_registers(2)(711));                                                         
                                                                                                                                     
        global_tmr_voter(1)(712)  <=    (tmr_registers(0)(712) and tmr_registers(1)(712)) or                                            
                            (tmr_registers(1)(712) and tmr_registers(2)(712)) or                                                       
                            (tmr_registers(0)(712) and tmr_registers(2)(712));                                                         
                                                                                                                                     
        global_tmr_voter(1)(713)  <=    (tmr_registers(0)(713) and tmr_registers(1)(713)) or                                            
                            (tmr_registers(1)(713) and tmr_registers(2)(713)) or                                                       
                            (tmr_registers(0)(713) and tmr_registers(2)(713));                                                         
                                                                                                                                     
        global_tmr_voter(1)(714)  <=    (tmr_registers(0)(714) and tmr_registers(1)(714)) or                                            
                            (tmr_registers(1)(714) and tmr_registers(2)(714)) or                                                       
                            (tmr_registers(0)(714) and tmr_registers(2)(714));                                                         
                                                                                                                                     
        global_tmr_voter(1)(715)  <=    (tmr_registers(0)(715) and tmr_registers(1)(715)) or                                            
                            (tmr_registers(1)(715) and tmr_registers(2)(715)) or                                                       
                            (tmr_registers(0)(715) and tmr_registers(2)(715));                                                         
                                                                                                                                     
        global_tmr_voter(1)(716)  <=    (tmr_registers(0)(716) and tmr_registers(1)(716)) or                                            
                            (tmr_registers(1)(716) and tmr_registers(2)(716)) or                                                       
                            (tmr_registers(0)(716) and tmr_registers(2)(716));                                                         
                                                                                                                                     
        global_tmr_voter(1)(717)  <=    (tmr_registers(0)(717) and tmr_registers(1)(717)) or                                            
                            (tmr_registers(1)(717) and tmr_registers(2)(717)) or                                                       
                            (tmr_registers(0)(717) and tmr_registers(2)(717));                                                         
                                                                                                                                     
        global_tmr_voter(1)(718)  <=    (tmr_registers(0)(718) and tmr_registers(1)(718)) or                                            
                            (tmr_registers(1)(718) and tmr_registers(2)(718)) or                                                       
                            (tmr_registers(0)(718) and tmr_registers(2)(718));                                                         
                                                                                                                                     
        global_tmr_voter(1)(719)  <=    (tmr_registers(0)(719) and tmr_registers(1)(719)) or                                            
                            (tmr_registers(1)(719) and tmr_registers(2)(719)) or                                                       
                            (tmr_registers(0)(719) and tmr_registers(2)(719));                                                         
                                                                                                                                     
        global_tmr_voter(1)(720)  <=    (tmr_registers(0)(720) and tmr_registers(1)(720)) or                                            
                            (tmr_registers(1)(720) and tmr_registers(2)(720)) or                                                       
                            (tmr_registers(0)(720) and tmr_registers(2)(720));                                                         
                                                                                                                                     
        global_tmr_voter(1)(721)  <=    (tmr_registers(0)(721) and tmr_registers(1)(721)) or                                            
                            (tmr_registers(1)(721) and tmr_registers(2)(721)) or                                                       
                            (tmr_registers(0)(721) and tmr_registers(2)(721));                                                         
                                                                                                                                     
        global_tmr_voter(1)(722)  <=    (tmr_registers(0)(722) and tmr_registers(1)(722)) or                                            
                            (tmr_registers(1)(722) and tmr_registers(2)(722)) or                                                       
                            (tmr_registers(0)(722) and tmr_registers(2)(722));                                                         
                                                                                                                                     
        global_tmr_voter(1)(723)  <=    (tmr_registers(0)(723) and tmr_registers(1)(723)) or                                            
                            (tmr_registers(1)(723) and tmr_registers(2)(723)) or                                                       
                            (tmr_registers(0)(723) and tmr_registers(2)(723));                                                         
                                                                                                                                     
        global_tmr_voter(1)(724)  <=    (tmr_registers(0)(724) and tmr_registers(1)(724)) or                                            
                            (tmr_registers(1)(724) and tmr_registers(2)(724)) or                                                       
                            (tmr_registers(0)(724) and tmr_registers(2)(724));                                                         
                                                                                                                                     
        global_tmr_voter(1)(725)  <=    (tmr_registers(0)(725) and tmr_registers(1)(725)) or                                            
                            (tmr_registers(1)(725) and tmr_registers(2)(725)) or                                                       
                            (tmr_registers(0)(725) and tmr_registers(2)(725));                                                         
                                                                                                                                     
        global_tmr_voter(1)(726)  <=    (tmr_registers(0)(726) and tmr_registers(1)(726)) or                                            
                            (tmr_registers(1)(726) and tmr_registers(2)(726)) or                                                       
                            (tmr_registers(0)(726) and tmr_registers(2)(726));                                                         
                                                                                                                                     
        global_tmr_voter(1)(727)  <=    (tmr_registers(0)(727) and tmr_registers(1)(727)) or                                            
                            (tmr_registers(1)(727) and tmr_registers(2)(727)) or                                                       
                            (tmr_registers(0)(727) and tmr_registers(2)(727));                                                         
                                                                                                                                     
        global_tmr_voter(1)(728)  <=    (tmr_registers(0)(728) and tmr_registers(1)(728)) or                                            
                            (tmr_registers(1)(728) and tmr_registers(2)(728)) or                                                       
                            (tmr_registers(0)(728) and tmr_registers(2)(728));                                                         
                                                                                                                                     
        global_tmr_voter(1)(729)  <=    (tmr_registers(0)(729) and tmr_registers(1)(729)) or                                            
                            (tmr_registers(1)(729) and tmr_registers(2)(729)) or                                                       
                            (tmr_registers(0)(729) and tmr_registers(2)(729));                                                         
                                                                                                                                     
        global_tmr_voter(1)(730)  <=    (tmr_registers(0)(730) and tmr_registers(1)(730)) or                                            
                            (tmr_registers(1)(730) and tmr_registers(2)(730)) or                                                       
                            (tmr_registers(0)(730) and tmr_registers(2)(730));                                                         
                                                                                                                                     
        global_tmr_voter(1)(731)  <=    (tmr_registers(0)(731) and tmr_registers(1)(731)) or                                            
                            (tmr_registers(1)(731) and tmr_registers(2)(731)) or                                                       
                            (tmr_registers(0)(731) and tmr_registers(2)(731));                                                         
                                                                                                                                     
        global_tmr_voter(1)(732)  <=    (tmr_registers(0)(732) and tmr_registers(1)(732)) or                                            
                            (tmr_registers(1)(732) and tmr_registers(2)(732)) or                                                       
                            (tmr_registers(0)(732) and tmr_registers(2)(732));                                                         
                                                                                                                                     
        global_tmr_voter(1)(733)  <=    (tmr_registers(0)(733) and tmr_registers(1)(733)) or                                            
                            (tmr_registers(1)(733) and tmr_registers(2)(733)) or                                                       
                            (tmr_registers(0)(733) and tmr_registers(2)(733));                                                         
                                                                                                                                     
        global_tmr_voter(1)(734)  <=    (tmr_registers(0)(734) and tmr_registers(1)(734)) or                                            
                            (tmr_registers(1)(734) and tmr_registers(2)(734)) or                                                       
                            (tmr_registers(0)(734) and tmr_registers(2)(734));                                                         
                                                                                                                                     
        global_tmr_voter(1)(735)  <=    (tmr_registers(0)(735) and tmr_registers(1)(735)) or                                            
                            (tmr_registers(1)(735) and tmr_registers(2)(735)) or                                                       
                            (tmr_registers(0)(735) and tmr_registers(2)(735));                                                         
                                                                                                                                     
        global_tmr_voter(1)(736)  <=    (tmr_registers(0)(736) and tmr_registers(1)(736)) or                                            
                            (tmr_registers(1)(736) and tmr_registers(2)(736)) or                                                       
                            (tmr_registers(0)(736) and tmr_registers(2)(736));                                                         
                                                                                                                                     
        global_tmr_voter(1)(737)  <=    (tmr_registers(0)(737) and tmr_registers(1)(737)) or                                            
                            (tmr_registers(1)(737) and tmr_registers(2)(737)) or                                                       
                            (tmr_registers(0)(737) and tmr_registers(2)(737));                                                         
                                                                                                                                     
        global_tmr_voter(1)(738)  <=    (tmr_registers(0)(738) and tmr_registers(1)(738)) or                                            
                            (tmr_registers(1)(738) and tmr_registers(2)(738)) or                                                       
                            (tmr_registers(0)(738) and tmr_registers(2)(738));                                                         
                                                                                                                                     
        global_tmr_voter(1)(739)  <=    (tmr_registers(0)(739) and tmr_registers(1)(739)) or                                            
                            (tmr_registers(1)(739) and tmr_registers(2)(739)) or                                                       
                            (tmr_registers(0)(739) and tmr_registers(2)(739));                                                         
                                                                                                                                     
        global_tmr_voter(1)(740)  <=    (tmr_registers(0)(740) and tmr_registers(1)(740)) or                                            
                            (tmr_registers(1)(740) and tmr_registers(2)(740)) or                                                       
                            (tmr_registers(0)(740) and tmr_registers(2)(740));                                                         
                                                                                                                                     
        global_tmr_voter(1)(741)  <=    (tmr_registers(0)(741) and tmr_registers(1)(741)) or                                            
                            (tmr_registers(1)(741) and tmr_registers(2)(741)) or                                                       
                            (tmr_registers(0)(741) and tmr_registers(2)(741));                                                         
                                                                                                                                     
        global_tmr_voter(1)(742)  <=    (tmr_registers(0)(742) and tmr_registers(1)(742)) or                                            
                            (tmr_registers(1)(742) and tmr_registers(2)(742)) or                                                       
                            (tmr_registers(0)(742) and tmr_registers(2)(742));                                                         
                                                                                                                                     
        global_tmr_voter(1)(743)  <=    (tmr_registers(0)(743) and tmr_registers(1)(743)) or                                            
                            (tmr_registers(1)(743) and tmr_registers(2)(743)) or                                                       
                            (tmr_registers(0)(743) and tmr_registers(2)(743));                                                         
                                                                                                                                     
        global_tmr_voter(1)(744)  <=    (tmr_registers(0)(744) and tmr_registers(1)(744)) or                                            
                            (tmr_registers(1)(744) and tmr_registers(2)(744)) or                                                       
                            (tmr_registers(0)(744) and tmr_registers(2)(744));                                                         
                                                                                                                                     
        global_tmr_voter(1)(745)  <=    (tmr_registers(0)(745) and tmr_registers(1)(745)) or                                            
                            (tmr_registers(1)(745) and tmr_registers(2)(745)) or                                                       
                            (tmr_registers(0)(745) and tmr_registers(2)(745));                                                         
                                                                                                                                     
        global_tmr_voter(1)(746)  <=    (tmr_registers(0)(746) and tmr_registers(1)(746)) or                                            
                            (tmr_registers(1)(746) and tmr_registers(2)(746)) or                                                       
                            (tmr_registers(0)(746) and tmr_registers(2)(746));                                                         
                                                                                                                                     
        global_tmr_voter(1)(747)  <=    (tmr_registers(0)(747) and tmr_registers(1)(747)) or                                            
                            (tmr_registers(1)(747) and tmr_registers(2)(747)) or                                                       
                            (tmr_registers(0)(747) and tmr_registers(2)(747));                                                         
                                                                                                                                     
        global_tmr_voter(1)(748)  <=    (tmr_registers(0)(748) and tmr_registers(1)(748)) or                                            
                            (tmr_registers(1)(748) and tmr_registers(2)(748)) or                                                       
                            (tmr_registers(0)(748) and tmr_registers(2)(748));                                                         
                                                                                                                                     
        global_tmr_voter(1)(749)  <=    (tmr_registers(0)(749) and tmr_registers(1)(749)) or                                            
                            (tmr_registers(1)(749) and tmr_registers(2)(749)) or                                                       
                            (tmr_registers(0)(749) and tmr_registers(2)(749));                                                         
                                                                                                                                     
        global_tmr_voter(1)(750)  <=    (tmr_registers(0)(750) and tmr_registers(1)(750)) or                                            
                            (tmr_registers(1)(750) and tmr_registers(2)(750)) or                                                       
                            (tmr_registers(0)(750) and tmr_registers(2)(750));                                                         
                                                                                                                                     
        global_tmr_voter(1)(751)  <=    (tmr_registers(0)(751) and tmr_registers(1)(751)) or                                            
                            (tmr_registers(1)(751) and tmr_registers(2)(751)) or                                                       
                            (tmr_registers(0)(751) and tmr_registers(2)(751));                                                         
                                                                                                                                     
        global_tmr_voter(1)(752)  <=    (tmr_registers(0)(752) and tmr_registers(1)(752)) or                                            
                            (tmr_registers(1)(752) and tmr_registers(2)(752)) or                                                       
                            (tmr_registers(0)(752) and tmr_registers(2)(752));                                                         
                                                                                                                                     
        global_tmr_voter(1)(753)  <=    (tmr_registers(0)(753) and tmr_registers(1)(753)) or                                            
                            (tmr_registers(1)(753) and tmr_registers(2)(753)) or                                                       
                            (tmr_registers(0)(753) and tmr_registers(2)(753));                                                         
                                                                                                                                     
        global_tmr_voter(1)(754)  <=    (tmr_registers(0)(754) and tmr_registers(1)(754)) or                                            
                            (tmr_registers(1)(754) and tmr_registers(2)(754)) or                                                       
                            (tmr_registers(0)(754) and tmr_registers(2)(754));                                                         
                                                                                                                                     
        global_tmr_voter(1)(755)  <=    (tmr_registers(0)(755) and tmr_registers(1)(755)) or                                            
                            (tmr_registers(1)(755) and tmr_registers(2)(755)) or                                                       
                            (tmr_registers(0)(755) and tmr_registers(2)(755));                                                         
                                                                                                                                     
        global_tmr_voter(1)(756)  <=    (tmr_registers(0)(756) and tmr_registers(1)(756)) or                                            
                            (tmr_registers(1)(756) and tmr_registers(2)(756)) or                                                       
                            (tmr_registers(0)(756) and tmr_registers(2)(756));                                                         
                                                                                                                                     
        global_tmr_voter(1)(757)  <=    (tmr_registers(0)(757) and tmr_registers(1)(757)) or                                            
                            (tmr_registers(1)(757) and tmr_registers(2)(757)) or                                                       
                            (tmr_registers(0)(757) and tmr_registers(2)(757));                                                         
                                                                                                                                     
        global_tmr_voter(1)(758)  <=    (tmr_registers(0)(758) and tmr_registers(1)(758)) or                                            
                            (tmr_registers(1)(758) and tmr_registers(2)(758)) or                                                       
                            (tmr_registers(0)(758) and tmr_registers(2)(758));                                                         
                                                                                                                                     
        global_tmr_voter(1)(759)  <=    (tmr_registers(0)(759) and tmr_registers(1)(759)) or                                            
                            (tmr_registers(1)(759) and tmr_registers(2)(759)) or                                                       
                            (tmr_registers(0)(759) and tmr_registers(2)(759));                                                         
                                                                                                                                     
        global_tmr_voter(1)(760)  <=    (tmr_registers(0)(760) and tmr_registers(1)(760)) or                                            
                            (tmr_registers(1)(760) and tmr_registers(2)(760)) or                                                       
                            (tmr_registers(0)(760) and tmr_registers(2)(760));                                                         
                                                                                                                                     
        global_tmr_voter(1)(761)  <=    (tmr_registers(0)(761) and tmr_registers(1)(761)) or                                            
                            (tmr_registers(1)(761) and tmr_registers(2)(761)) or                                                       
                            (tmr_registers(0)(761) and tmr_registers(2)(761));                                                         
                                                                                                                                     
        global_tmr_voter(1)(762)  <=    (tmr_registers(0)(762) and tmr_registers(1)(762)) or                                            
                            (tmr_registers(1)(762) and tmr_registers(2)(762)) or                                                       
                            (tmr_registers(0)(762) and tmr_registers(2)(762));                                                         
                                                                                                                                     
        global_tmr_voter(1)(763)  <=    (tmr_registers(0)(763) and tmr_registers(1)(763)) or                                            
                            (tmr_registers(1)(763) and tmr_registers(2)(763)) or                                                       
                            (tmr_registers(0)(763) and tmr_registers(2)(763));                                                         
                                                                                                                                     
        global_tmr_voter(1)(764)  <=    (tmr_registers(0)(764) and tmr_registers(1)(764)) or                                            
                            (tmr_registers(1)(764) and tmr_registers(2)(764)) or                                                       
                            (tmr_registers(0)(764) and tmr_registers(2)(764));                                                         
                                                                                                                                     
        global_tmr_voter(1)(765)  <=    (tmr_registers(0)(765) and tmr_registers(1)(765)) or                                            
                            (tmr_registers(1)(765) and tmr_registers(2)(765)) or                                                       
                            (tmr_registers(0)(765) and tmr_registers(2)(765));                                                         
                                                                                                                                     
        global_tmr_voter(1)(766)  <=    (tmr_registers(0)(766) and tmr_registers(1)(766)) or                                            
                            (tmr_registers(1)(766) and tmr_registers(2)(766)) or                                                       
                            (tmr_registers(0)(766) and tmr_registers(2)(766));                                                         
                                                                                                                                     
        global_tmr_voter(1)(767)  <=    (tmr_registers(0)(767) and tmr_registers(1)(767)) or                                            
                            (tmr_registers(1)(767) and tmr_registers(2)(767)) or                                                       
                            (tmr_registers(0)(767) and tmr_registers(2)(767));                                                         
                                                                                                                                     
        global_tmr_voter(1)(768)  <=    (tmr_registers(0)(768) and tmr_registers(1)(768)) or                                            
                            (tmr_registers(1)(768) and tmr_registers(2)(768)) or                                                       
                            (tmr_registers(0)(768) and tmr_registers(2)(768));                                                         
                                                                                                                                     
        global_tmr_voter(1)(769)  <=    (tmr_registers(0)(769) and tmr_registers(1)(769)) or                                            
                            (tmr_registers(1)(769) and tmr_registers(2)(769)) or                                                       
                            (tmr_registers(0)(769) and tmr_registers(2)(769));                                                         
                                                                                                                                     
        global_tmr_voter(1)(770)  <=    (tmr_registers(0)(770) and tmr_registers(1)(770)) or                                            
                            (tmr_registers(1)(770) and tmr_registers(2)(770)) or                                                       
                            (tmr_registers(0)(770) and tmr_registers(2)(770));                                                         
                                                                                                                                     
        global_tmr_voter(1)(771)  <=    (tmr_registers(0)(771) and tmr_registers(1)(771)) or                                            
                            (tmr_registers(1)(771) and tmr_registers(2)(771)) or                                                       
                            (tmr_registers(0)(771) and tmr_registers(2)(771));                                                         
                                                                                                                                     
        global_tmr_voter(1)(772)  <=    (tmr_registers(0)(772) and tmr_registers(1)(772)) or                                            
                            (tmr_registers(1)(772) and tmr_registers(2)(772)) or                                                       
                            (tmr_registers(0)(772) and tmr_registers(2)(772));                                                         
                                                                                                                                     
        global_tmr_voter(1)(773)  <=    (tmr_registers(0)(773) and tmr_registers(1)(773)) or                                            
                            (tmr_registers(1)(773) and tmr_registers(2)(773)) or                                                       
                            (tmr_registers(0)(773) and tmr_registers(2)(773));                                                         
                                                                                                                                     
        global_tmr_voter(1)(774)  <=    (tmr_registers(0)(774) and tmr_registers(1)(774)) or                                            
                            (tmr_registers(1)(774) and tmr_registers(2)(774)) or                                                       
                            (tmr_registers(0)(774) and tmr_registers(2)(774));                                                         
                                                                                                                                     
        global_tmr_voter(1)(775)  <=    (tmr_registers(0)(775) and tmr_registers(1)(775)) or                                            
                            (tmr_registers(1)(775) and tmr_registers(2)(775)) or                                                       
                            (tmr_registers(0)(775) and tmr_registers(2)(775));                                                         
                                                                                                                                     
        global_tmr_voter(1)(776)  <=    (tmr_registers(0)(776) and tmr_registers(1)(776)) or                                            
                            (tmr_registers(1)(776) and tmr_registers(2)(776)) or                                                       
                            (tmr_registers(0)(776) and tmr_registers(2)(776));                                                         
                                                                                                                                     
        global_tmr_voter(1)(777)  <=    (tmr_registers(0)(777) and tmr_registers(1)(777)) or                                            
                            (tmr_registers(1)(777) and tmr_registers(2)(777)) or                                                       
                            (tmr_registers(0)(777) and tmr_registers(2)(777));                                                         
                                                                                                                                     
        global_tmr_voter(1)(778)  <=    (tmr_registers(0)(778) and tmr_registers(1)(778)) or                                            
                            (tmr_registers(1)(778) and tmr_registers(2)(778)) or                                                       
                            (tmr_registers(0)(778) and tmr_registers(2)(778));                                                         
                                                                                                                                     
        global_tmr_voter(1)(779)  <=    (tmr_registers(0)(779) and tmr_registers(1)(779)) or                                            
                            (tmr_registers(1)(779) and tmr_registers(2)(779)) or                                                       
                            (tmr_registers(0)(779) and tmr_registers(2)(779));                                                         
                                                                                                                                     
        global_tmr_voter(1)(780)  <=    (tmr_registers(0)(780) and tmr_registers(1)(780)) or                                            
                            (tmr_registers(1)(780) and tmr_registers(2)(780)) or                                                       
                            (tmr_registers(0)(780) and tmr_registers(2)(780));                                                         
                                                                                                                                     
        global_tmr_voter(1)(781)  <=    (tmr_registers(0)(781) and tmr_registers(1)(781)) or                                            
                            (tmr_registers(1)(781) and tmr_registers(2)(781)) or                                                       
                            (tmr_registers(0)(781) and tmr_registers(2)(781));                                                         
                                                                                                                                     
        global_tmr_voter(1)(782)  <=    (tmr_registers(0)(782) and tmr_registers(1)(782)) or                                            
                            (tmr_registers(1)(782) and tmr_registers(2)(782)) or                                                       
                            (tmr_registers(0)(782) and tmr_registers(2)(782));                                                         
                                                                                                                                     
        global_tmr_voter(1)(783)  <=    (tmr_registers(0)(783) and tmr_registers(1)(783)) or                                            
                            (tmr_registers(1)(783) and tmr_registers(2)(783)) or                                                       
                            (tmr_registers(0)(783) and tmr_registers(2)(783));                                                         
                                                                                                                                     
        global_tmr_voter(1)(784)  <=    (tmr_registers(0)(784) and tmr_registers(1)(784)) or                                            
                            (tmr_registers(1)(784) and tmr_registers(2)(784)) or                                                       
                            (tmr_registers(0)(784) and tmr_registers(2)(784));                                                         
                                                                                                                                     
        global_tmr_voter(1)(785)  <=    (tmr_registers(0)(785) and tmr_registers(1)(785)) or                                            
                            (tmr_registers(1)(785) and tmr_registers(2)(785)) or                                                       
                            (tmr_registers(0)(785) and tmr_registers(2)(785));                                                         
                                                                                                                                     
        global_tmr_voter(1)(786)  <=    (tmr_registers(0)(786) and tmr_registers(1)(786)) or                                            
                            (tmr_registers(1)(786) and tmr_registers(2)(786)) or                                                       
                            (tmr_registers(0)(786) and tmr_registers(2)(786));                                                         
                                                                                                                                     
        global_tmr_voter(1)(787)  <=    (tmr_registers(0)(787) and tmr_registers(1)(787)) or                                            
                            (tmr_registers(1)(787) and tmr_registers(2)(787)) or                                                       
                            (tmr_registers(0)(787) and tmr_registers(2)(787));                                                         
                                                                                                                                     
        global_tmr_voter(1)(788)  <=    (tmr_registers(0)(788) and tmr_registers(1)(788)) or                                            
                            (tmr_registers(1)(788) and tmr_registers(2)(788)) or                                                       
                            (tmr_registers(0)(788) and tmr_registers(2)(788));                                                         
                                                                                                                                     
        global_tmr_voter(1)(789)  <=    (tmr_registers(0)(789) and tmr_registers(1)(789)) or                                            
                            (tmr_registers(1)(789) and tmr_registers(2)(789)) or                                                       
                            (tmr_registers(0)(789) and tmr_registers(2)(789));                                                         
                                                                                                                                     
        global_tmr_voter(1)(790)  <=    (tmr_registers(0)(790) and tmr_registers(1)(790)) or                                            
                            (tmr_registers(1)(790) and tmr_registers(2)(790)) or                                                       
                            (tmr_registers(0)(790) and tmr_registers(2)(790));                                                         
                                                                                                                                     
        global_tmr_voter(1)(791)  <=    (tmr_registers(0)(791) and tmr_registers(1)(791)) or                                            
                            (tmr_registers(1)(791) and tmr_registers(2)(791)) or                                                       
                            (tmr_registers(0)(791) and tmr_registers(2)(791));                                                         
                                                                                                                                     
        global_tmr_voter(1)(792)  <=    (tmr_registers(0)(792) and tmr_registers(1)(792)) or                                            
                            (tmr_registers(1)(792) and tmr_registers(2)(792)) or                                                       
                            (tmr_registers(0)(792) and tmr_registers(2)(792));                                                         
                                                                                                                                     
        global_tmr_voter(1)(793)  <=    (tmr_registers(0)(793) and tmr_registers(1)(793)) or                                            
                            (tmr_registers(1)(793) and tmr_registers(2)(793)) or                                                       
                            (tmr_registers(0)(793) and tmr_registers(2)(793));                                                         
                                                                                                                                     
        global_tmr_voter(1)(794)  <=    (tmr_registers(0)(794) and tmr_registers(1)(794)) or                                            
                            (tmr_registers(1)(794) and tmr_registers(2)(794)) or                                                       
                            (tmr_registers(0)(794) and tmr_registers(2)(794));                                                         
                                                                                                                                     
        global_tmr_voter(1)(795)  <=    (tmr_registers(0)(795) and tmr_registers(1)(795)) or                                            
                            (tmr_registers(1)(795) and tmr_registers(2)(795)) or                                                       
                            (tmr_registers(0)(795) and tmr_registers(2)(795));                                                         
                                                                                                                                     
        global_tmr_voter(1)(796)  <=    (tmr_registers(0)(796) and tmr_registers(1)(796)) or                                            
                            (tmr_registers(1)(796) and tmr_registers(2)(796)) or                                                       
                            (tmr_registers(0)(796) and tmr_registers(2)(796));                                                         
                                                                                                                                     
        global_tmr_voter(1)(797)  <=    (tmr_registers(0)(797) and tmr_registers(1)(797)) or                                            
                            (tmr_registers(1)(797) and tmr_registers(2)(797)) or                                                       
                            (tmr_registers(0)(797) and tmr_registers(2)(797));                                                         
                                                                                                                                     
        global_tmr_voter(1)(798)  <=    (tmr_registers(0)(798) and tmr_registers(1)(798)) or                                            
                            (tmr_registers(1)(798) and tmr_registers(2)(798)) or                                                       
                            (tmr_registers(0)(798) and tmr_registers(2)(798));                                                         
                                                                                                                                     
        global_tmr_voter(1)(799)  <=    (tmr_registers(0)(799) and tmr_registers(1)(799)) or                                            
                            (tmr_registers(1)(799) and tmr_registers(2)(799)) or                                                       
                            (tmr_registers(0)(799) and tmr_registers(2)(799));                                                         
                                                                                                                                     
        global_tmr_voter(1)(800)  <=    (tmr_registers(0)(800) and tmr_registers(1)(800)) or                                            
                            (tmr_registers(1)(800) and tmr_registers(2)(800)) or                                                       
                            (tmr_registers(0)(800) and tmr_registers(2)(800));                                                         
                                                                                                                                     
        global_tmr_voter(1)(801)  <=    (tmr_registers(0)(801) and tmr_registers(1)(801)) or                                            
                            (tmr_registers(1)(801) and tmr_registers(2)(801)) or                                                       
                            (tmr_registers(0)(801) and tmr_registers(2)(801));                                                         
                                                                                                                                     
        global_tmr_voter(1)(802)  <=    (tmr_registers(0)(802) and tmr_registers(1)(802)) or                                            
                            (tmr_registers(1)(802) and tmr_registers(2)(802)) or                                                       
                            (tmr_registers(0)(802) and tmr_registers(2)(802));                                                         
                                                                                                                                     
        global_tmr_voter(1)(803)  <=    (tmr_registers(0)(803) and tmr_registers(1)(803)) or                                            
                            (tmr_registers(1)(803) and tmr_registers(2)(803)) or                                                       
                            (tmr_registers(0)(803) and tmr_registers(2)(803));                                                         
                                                                                                                                     
        global_tmr_voter(1)(804)  <=    (tmr_registers(0)(804) and tmr_registers(1)(804)) or                                            
                            (tmr_registers(1)(804) and tmr_registers(2)(804)) or                                                       
                            (tmr_registers(0)(804) and tmr_registers(2)(804));                                                         
                                                                                                                                     
        global_tmr_voter(1)(805)  <=    (tmr_registers(0)(805) and tmr_registers(1)(805)) or                                            
                            (tmr_registers(1)(805) and tmr_registers(2)(805)) or                                                       
                            (tmr_registers(0)(805) and tmr_registers(2)(805));                                                         
                                                                                                                                     
        global_tmr_voter(1)(806)  <=    (tmr_registers(0)(806) and tmr_registers(1)(806)) or                                            
                            (tmr_registers(1)(806) and tmr_registers(2)(806)) or                                                       
                            (tmr_registers(0)(806) and tmr_registers(2)(806));                                                         
                                                                                                                                     
        global_tmr_voter(1)(807)  <=    (tmr_registers(0)(807) and tmr_registers(1)(807)) or                                            
                            (tmr_registers(1)(807) and tmr_registers(2)(807)) or                                                       
                            (tmr_registers(0)(807) and tmr_registers(2)(807));                                                         
                                                                                                                                     
        global_tmr_voter(1)(808)  <=    (tmr_registers(0)(808) and tmr_registers(1)(808)) or                                            
                            (tmr_registers(1)(808) and tmr_registers(2)(808)) or                                                       
                            (tmr_registers(0)(808) and tmr_registers(2)(808));                                                         
                                                                                                                                     
        global_tmr_voter(1)(809)  <=    (tmr_registers(0)(809) and tmr_registers(1)(809)) or                                            
                            (tmr_registers(1)(809) and tmr_registers(2)(809)) or                                                       
                            (tmr_registers(0)(809) and tmr_registers(2)(809));                                                         
                                                                                                                                     
        global_tmr_voter(1)(810)  <=    (tmr_registers(0)(810) and tmr_registers(1)(810)) or                                            
                            (tmr_registers(1)(810) and tmr_registers(2)(810)) or                                                       
                            (tmr_registers(0)(810) and tmr_registers(2)(810));                                                         
                                                                                                                                     
        global_tmr_voter(1)(811)  <=    (tmr_registers(0)(811) and tmr_registers(1)(811)) or                                            
                            (tmr_registers(1)(811) and tmr_registers(2)(811)) or                                                       
                            (tmr_registers(0)(811) and tmr_registers(2)(811));                                                         
                                                                                                                                     
        global_tmr_voter(1)(812)  <=    (tmr_registers(0)(812) and tmr_registers(1)(812)) or                                            
                            (tmr_registers(1)(812) and tmr_registers(2)(812)) or                                                       
                            (tmr_registers(0)(812) and tmr_registers(2)(812));                                                         
                                                                                                                                     
        global_tmr_voter(1)(813)  <=    (tmr_registers(0)(813) and tmr_registers(1)(813)) or                                            
                            (tmr_registers(1)(813) and tmr_registers(2)(813)) or                                                       
                            (tmr_registers(0)(813) and tmr_registers(2)(813));                                                         
                                                                                                                                     
        global_tmr_voter(1)(814)  <=    (tmr_registers(0)(814) and tmr_registers(1)(814)) or                                            
                            (tmr_registers(1)(814) and tmr_registers(2)(814)) or                                                       
                            (tmr_registers(0)(814) and tmr_registers(2)(814));                                                         
                                                                                                                                     
        global_tmr_voter(1)(815)  <=    (tmr_registers(0)(815) and tmr_registers(1)(815)) or                                            
                            (tmr_registers(1)(815) and tmr_registers(2)(815)) or                                                       
                            (tmr_registers(0)(815) and tmr_registers(2)(815));                                                         
                                                                                                                                     
        global_tmr_voter(1)(816)  <=    (tmr_registers(0)(816) and tmr_registers(1)(816)) or                                            
                            (tmr_registers(1)(816) and tmr_registers(2)(816)) or                                                       
                            (tmr_registers(0)(816) and tmr_registers(2)(816));                                                         
                                                                                                                                     
        global_tmr_voter(1)(817)  <=    (tmr_registers(0)(817) and tmr_registers(1)(817)) or                                            
                            (tmr_registers(1)(817) and tmr_registers(2)(817)) or                                                       
                            (tmr_registers(0)(817) and tmr_registers(2)(817));                                                         
                                                                                                                                     
        global_tmr_voter(1)(818)  <=    (tmr_registers(0)(818) and tmr_registers(1)(818)) or                                            
                            (tmr_registers(1)(818) and tmr_registers(2)(818)) or                                                       
                            (tmr_registers(0)(818) and tmr_registers(2)(818));                                                         
                                                                                                                                     
        global_tmr_voter(1)(819)  <=    (tmr_registers(0)(819) and tmr_registers(1)(819)) or                                            
                            (tmr_registers(1)(819) and tmr_registers(2)(819)) or                                                       
                            (tmr_registers(0)(819) and tmr_registers(2)(819));                                                         
                                                                                                                                     
        global_tmr_voter(1)(820)  <=    (tmr_registers(0)(820) and tmr_registers(1)(820)) or                                            
                            (tmr_registers(1)(820) and tmr_registers(2)(820)) or                                                       
                            (tmr_registers(0)(820) and tmr_registers(2)(820));                                                         
                                                                                                                                     
        global_tmr_voter(1)(821)  <=    (tmr_registers(0)(821) and tmr_registers(1)(821)) or                                            
                            (tmr_registers(1)(821) and tmr_registers(2)(821)) or                                                       
                            (tmr_registers(0)(821) and tmr_registers(2)(821));                                                         
                                                                                                                                     
        global_tmr_voter(1)(822)  <=    (tmr_registers(0)(822) and tmr_registers(1)(822)) or                                            
                            (tmr_registers(1)(822) and tmr_registers(2)(822)) or                                                       
                            (tmr_registers(0)(822) and tmr_registers(2)(822));                                                         
                                                                                                                                     
        global_tmr_voter(1)(823)  <=    (tmr_registers(0)(823) and tmr_registers(1)(823)) or                                            
                            (tmr_registers(1)(823) and tmr_registers(2)(823)) or                                                       
                            (tmr_registers(0)(823) and tmr_registers(2)(823));                                                         
                                                                                                                                     
        global_tmr_voter(1)(824)  <=    (tmr_registers(0)(824) and tmr_registers(1)(824)) or                                            
                            (tmr_registers(1)(824) and tmr_registers(2)(824)) or                                                       
                            (tmr_registers(0)(824) and tmr_registers(2)(824));                                                         
                                                                                                                                     
        global_tmr_voter(1)(825)  <=    (tmr_registers(0)(825) and tmr_registers(1)(825)) or                                            
                            (tmr_registers(1)(825) and tmr_registers(2)(825)) or                                                       
                            (tmr_registers(0)(825) and tmr_registers(2)(825));                                                         
                                                                                                                                     
        global_tmr_voter(1)(826)  <=    (tmr_registers(0)(826) and tmr_registers(1)(826)) or                                            
                            (tmr_registers(1)(826) and tmr_registers(2)(826)) or                                                       
                            (tmr_registers(0)(826) and tmr_registers(2)(826));                                                         
                                                                                                                                     
        global_tmr_voter(1)(827)  <=    (tmr_registers(0)(827) and tmr_registers(1)(827)) or                                            
                            (tmr_registers(1)(827) and tmr_registers(2)(827)) or                                                       
                            (tmr_registers(0)(827) and tmr_registers(2)(827));                                                         
                                                                                                                                     
        global_tmr_voter(1)(828)  <=    (tmr_registers(0)(828) and tmr_registers(1)(828)) or                                            
                            (tmr_registers(1)(828) and tmr_registers(2)(828)) or                                                       
                            (tmr_registers(0)(828) and tmr_registers(2)(828));                                                         
                                                                                                                                     
        global_tmr_voter(1)(829)  <=    (tmr_registers(0)(829) and tmr_registers(1)(829)) or                                            
                            (tmr_registers(1)(829) and tmr_registers(2)(829)) or                                                       
                            (tmr_registers(0)(829) and tmr_registers(2)(829));                                                         
                                                                                                                                     
        global_tmr_voter(1)(830)  <=    (tmr_registers(0)(830) and tmr_registers(1)(830)) or                                            
                            (tmr_registers(1)(830) and tmr_registers(2)(830)) or                                                       
                            (tmr_registers(0)(830) and tmr_registers(2)(830));                                                         
                                                                                                                                     
        global_tmr_voter(1)(831)  <=    (tmr_registers(0)(831) and tmr_registers(1)(831)) or                                            
                            (tmr_registers(1)(831) and tmr_registers(2)(831)) or                                                       
                            (tmr_registers(0)(831) and tmr_registers(2)(831));                                                         
                                                                                                                                     
        global_tmr_voter(1)(832)  <=    (tmr_registers(0)(832) and tmr_registers(1)(832)) or                                            
                            (tmr_registers(1)(832) and tmr_registers(2)(832)) or                                                       
                            (tmr_registers(0)(832) and tmr_registers(2)(832));                                                         
                                                                                                                                     
        global_tmr_voter(1)(833)  <=    (tmr_registers(0)(833) and tmr_registers(1)(833)) or                                            
                            (tmr_registers(1)(833) and tmr_registers(2)(833)) or                                                       
                            (tmr_registers(0)(833) and tmr_registers(2)(833));                                                         
                                                                                                                                     
        global_tmr_voter(1)(834)  <=    (tmr_registers(0)(834) and tmr_registers(1)(834)) or                                            
                            (tmr_registers(1)(834) and tmr_registers(2)(834)) or                                                       
                            (tmr_registers(0)(834) and tmr_registers(2)(834));                                                         
                                                                                                                                     
        global_tmr_voter(1)(835)  <=    (tmr_registers(0)(835) and tmr_registers(1)(835)) or                                            
                            (tmr_registers(1)(835) and tmr_registers(2)(835)) or                                                       
                            (tmr_registers(0)(835) and tmr_registers(2)(835));                                                         
                                                                                                                                     
        global_tmr_voter(1)(836)  <=    (tmr_registers(0)(836) and tmr_registers(1)(836)) or                                            
                            (tmr_registers(1)(836) and tmr_registers(2)(836)) or                                                       
                            (tmr_registers(0)(836) and tmr_registers(2)(836));                                                         
                                                                                                                                     
        global_tmr_voter(1)(837)  <=    (tmr_registers(0)(837) and tmr_registers(1)(837)) or                                            
                            (tmr_registers(1)(837) and tmr_registers(2)(837)) or                                                       
                            (tmr_registers(0)(837) and tmr_registers(2)(837));                                                         
                                                                                                                                     
        global_tmr_voter(1)(838)  <=    (tmr_registers(0)(838) and tmr_registers(1)(838)) or                                            
                            (tmr_registers(1)(838) and tmr_registers(2)(838)) or                                                       
                            (tmr_registers(0)(838) and tmr_registers(2)(838));                                                         
                                                                                                                                     
        global_tmr_voter(1)(839)  <=    (tmr_registers(0)(839) and tmr_registers(1)(839)) or                                            
                            (tmr_registers(1)(839) and tmr_registers(2)(839)) or                                                       
                            (tmr_registers(0)(839) and tmr_registers(2)(839));                                                         
                                                                                                                                     
        global_tmr_voter(1)(840)  <=    (tmr_registers(0)(840) and tmr_registers(1)(840)) or                                            
                            (tmr_registers(1)(840) and tmr_registers(2)(840)) or                                                       
                            (tmr_registers(0)(840) and tmr_registers(2)(840));                                                         
                                                                                                                                     
        global_tmr_voter(1)(841)  <=    (tmr_registers(0)(841) and tmr_registers(1)(841)) or                                            
                            (tmr_registers(1)(841) and tmr_registers(2)(841)) or                                                       
                            (tmr_registers(0)(841) and tmr_registers(2)(841));                                                         
                                                                                                                                     
        global_tmr_voter(1)(842)  <=    (tmr_registers(0)(842) and tmr_registers(1)(842)) or                                            
                            (tmr_registers(1)(842) and tmr_registers(2)(842)) or                                                       
                            (tmr_registers(0)(842) and tmr_registers(2)(842));                                                         
                                                                                                                                     
        global_tmr_voter(1)(843)  <=    (tmr_registers(0)(843) and tmr_registers(1)(843)) or                                            
                            (tmr_registers(1)(843) and tmr_registers(2)(843)) or                                                       
                            (tmr_registers(0)(843) and tmr_registers(2)(843));                                                         
                                                                                                                                     
        global_tmr_voter(1)(844)  <=    (tmr_registers(0)(844) and tmr_registers(1)(844)) or                                            
                            (tmr_registers(1)(844) and tmr_registers(2)(844)) or                                                       
                            (tmr_registers(0)(844) and tmr_registers(2)(844));                                                         
                                                                                                                                     
        global_tmr_voter(1)(845)  <=    (tmr_registers(0)(845) and tmr_registers(1)(845)) or                                            
                            (tmr_registers(1)(845) and tmr_registers(2)(845)) or                                                       
                            (tmr_registers(0)(845) and tmr_registers(2)(845));                                                         
                                                                                                                                     
        global_tmr_voter(1)(846)  <=    (tmr_registers(0)(846) and tmr_registers(1)(846)) or                                            
                            (tmr_registers(1)(846) and tmr_registers(2)(846)) or                                                       
                            (tmr_registers(0)(846) and tmr_registers(2)(846));                                                         
                                                                                                                                     
        global_tmr_voter(1)(847)  <=    (tmr_registers(0)(847) and tmr_registers(1)(847)) or                                            
                            (tmr_registers(1)(847) and tmr_registers(2)(847)) or                                                       
                            (tmr_registers(0)(847) and tmr_registers(2)(847));                                                         
                                                                                                                                     
        global_tmr_voter(1)(848)  <=    (tmr_registers(0)(848) and tmr_registers(1)(848)) or                                            
                            (tmr_registers(1)(848) and tmr_registers(2)(848)) or                                                       
                            (tmr_registers(0)(848) and tmr_registers(2)(848));                                                         
                                                                                                                                     
        global_tmr_voter(1)(849)  <=    (tmr_registers(0)(849) and tmr_registers(1)(849)) or                                            
                            (tmr_registers(1)(849) and tmr_registers(2)(849)) or                                                       
                            (tmr_registers(0)(849) and tmr_registers(2)(849));                                                         
                                                                                                                                     
        global_tmr_voter(1)(850)  <=    (tmr_registers(0)(850) and tmr_registers(1)(850)) or                                            
                            (tmr_registers(1)(850) and tmr_registers(2)(850)) or                                                       
                            (tmr_registers(0)(850) and tmr_registers(2)(850));                                                         
                                                                                                                                     
        global_tmr_voter(1)(851)  <=    (tmr_registers(0)(851) and tmr_registers(1)(851)) or                                            
                            (tmr_registers(1)(851) and tmr_registers(2)(851)) or                                                       
                            (tmr_registers(0)(851) and tmr_registers(2)(851));                                                         
                                                                                                                                     
        global_tmr_voter(1)(852)  <=    (tmr_registers(0)(852) and tmr_registers(1)(852)) or                                            
                            (tmr_registers(1)(852) and tmr_registers(2)(852)) or                                                       
                            (tmr_registers(0)(852) and tmr_registers(2)(852));                                                         
                                                                                                                                     
        global_tmr_voter(1)(853)  <=    (tmr_registers(0)(853) and tmr_registers(1)(853)) or                                            
                            (tmr_registers(1)(853) and tmr_registers(2)(853)) or                                                       
                            (tmr_registers(0)(853) and tmr_registers(2)(853));                                                         
                                                                                                                                     
        global_tmr_voter(1)(854)  <=    (tmr_registers(0)(854) and tmr_registers(1)(854)) or                                            
                            (tmr_registers(1)(854) and tmr_registers(2)(854)) or                                                       
                            (tmr_registers(0)(854) and tmr_registers(2)(854));                                                         
                                                                                                                                     
        global_tmr_voter(1)(855)  <=    (tmr_registers(0)(855) and tmr_registers(1)(855)) or                                            
                            (tmr_registers(1)(855) and tmr_registers(2)(855)) or                                                       
                            (tmr_registers(0)(855) and tmr_registers(2)(855));                                                         
                                                                                                                                     
        global_tmr_voter(1)(856)  <=    (tmr_registers(0)(856) and tmr_registers(1)(856)) or                                            
                            (tmr_registers(1)(856) and tmr_registers(2)(856)) or                                                       
                            (tmr_registers(0)(856) and tmr_registers(2)(856));                                                         
                                                                                                                                     
        global_tmr_voter(1)(857)  <=    (tmr_registers(0)(857) and tmr_registers(1)(857)) or                                            
                            (tmr_registers(1)(857) and tmr_registers(2)(857)) or                                                       
                            (tmr_registers(0)(857) and tmr_registers(2)(857));                                                         
                                                                                                                                     
        global_tmr_voter(1)(858)  <=    (tmr_registers(0)(858) and tmr_registers(1)(858)) or                                            
                            (tmr_registers(1)(858) and tmr_registers(2)(858)) or                                                       
                            (tmr_registers(0)(858) and tmr_registers(2)(858));                                                         
                                                                                                                                     
        global_tmr_voter(1)(859)  <=    (tmr_registers(0)(859) and tmr_registers(1)(859)) or                                            
                            (tmr_registers(1)(859) and tmr_registers(2)(859)) or                                                       
                            (tmr_registers(0)(859) and tmr_registers(2)(859));                                                         
                                                                                                                                     
        global_tmr_voter(1)(860)  <=    (tmr_registers(0)(860) and tmr_registers(1)(860)) or                                            
                            (tmr_registers(1)(860) and tmr_registers(2)(860)) or                                                       
                            (tmr_registers(0)(860) and tmr_registers(2)(860));                                                         
                                                                                                                                     
        global_tmr_voter(1)(861)  <=    (tmr_registers(0)(861) and tmr_registers(1)(861)) or                                            
                            (tmr_registers(1)(861) and tmr_registers(2)(861)) or                                                       
                            (tmr_registers(0)(861) and tmr_registers(2)(861));                                                         
                                                                                                                                     
        global_tmr_voter(1)(862)  <=    (tmr_registers(0)(862) and tmr_registers(1)(862)) or                                            
                            (tmr_registers(1)(862) and tmr_registers(2)(862)) or                                                       
                            (tmr_registers(0)(862) and tmr_registers(2)(862));                                                         
                                                                                                                                     
        global_tmr_voter(1)(863)  <=    (tmr_registers(0)(863) and tmr_registers(1)(863)) or                                            
                            (tmr_registers(1)(863) and tmr_registers(2)(863)) or                                                       
                            (tmr_registers(0)(863) and tmr_registers(2)(863));                                                         
                                                                                                                                     
        global_tmr_voter(1)(864)  <=    (tmr_registers(0)(864) and tmr_registers(1)(864)) or                                            
                            (tmr_registers(1)(864) and tmr_registers(2)(864)) or                                                       
                            (tmr_registers(0)(864) and tmr_registers(2)(864));                                                         
                                                                                                                                     
        global_tmr_voter(1)(865)  <=    (tmr_registers(0)(865) and tmr_registers(1)(865)) or                                            
                            (tmr_registers(1)(865) and tmr_registers(2)(865)) or                                                       
                            (tmr_registers(0)(865) and tmr_registers(2)(865));                                                         
                                                                                                                                     
        global_tmr_voter(1)(866)  <=    (tmr_registers(0)(866) and tmr_registers(1)(866)) or                                            
                            (tmr_registers(1)(866) and tmr_registers(2)(866)) or                                                       
                            (tmr_registers(0)(866) and tmr_registers(2)(866));                                                         
                                                                                                                                     
        global_tmr_voter(1)(867)  <=    (tmr_registers(0)(867) and tmr_registers(1)(867)) or                                            
                            (tmr_registers(1)(867) and tmr_registers(2)(867)) or                                                       
                            (tmr_registers(0)(867) and tmr_registers(2)(867));                                                         
                                                                                                                                     
        global_tmr_voter(1)(868)  <=    (tmr_registers(0)(868) and tmr_registers(1)(868)) or                                            
                            (tmr_registers(1)(868) and tmr_registers(2)(868)) or                                                       
                            (tmr_registers(0)(868) and tmr_registers(2)(868));                                                         
                                                                                                                                     
        global_tmr_voter(1)(869)  <=    (tmr_registers(0)(869) and tmr_registers(1)(869)) or                                            
                            (tmr_registers(1)(869) and tmr_registers(2)(869)) or                                                       
                            (tmr_registers(0)(869) and tmr_registers(2)(869));                                                         
                                                                                                                                     
        global_tmr_voter(1)(870)  <=    (tmr_registers(0)(870) and tmr_registers(1)(870)) or                                            
                            (tmr_registers(1)(870) and tmr_registers(2)(870)) or                                                       
                            (tmr_registers(0)(870) and tmr_registers(2)(870));                                                         
                                                                                                                                     
        global_tmr_voter(1)(871)  <=    (tmr_registers(0)(871) and tmr_registers(1)(871)) or                                            
                            (tmr_registers(1)(871) and tmr_registers(2)(871)) or                                                       
                            (tmr_registers(0)(871) and tmr_registers(2)(871));                                                         
                                                                                                                                     
        global_tmr_voter(1)(872)  <=    (tmr_registers(0)(872) and tmr_registers(1)(872)) or                                            
                            (tmr_registers(1)(872) and tmr_registers(2)(872)) or                                                       
                            (tmr_registers(0)(872) and tmr_registers(2)(872));                                                         
                                                                                                                                     
        global_tmr_voter(1)(873)  <=    (tmr_registers(0)(873) and tmr_registers(1)(873)) or                                            
                            (tmr_registers(1)(873) and tmr_registers(2)(873)) or                                                       
                            (tmr_registers(0)(873) and tmr_registers(2)(873));                                                         
                                                                                                                                     
        global_tmr_voter(1)(874)  <=    (tmr_registers(0)(874) and tmr_registers(1)(874)) or                                            
                            (tmr_registers(1)(874) and tmr_registers(2)(874)) or                                                       
                            (tmr_registers(0)(874) and tmr_registers(2)(874));                                                         
                                                                                                                                     
        global_tmr_voter(1)(875)  <=    (tmr_registers(0)(875) and tmr_registers(1)(875)) or                                            
                            (tmr_registers(1)(875) and tmr_registers(2)(875)) or                                                       
                            (tmr_registers(0)(875) and tmr_registers(2)(875));                                                         
                                                                                                                                     
        global_tmr_voter(1)(876)  <=    (tmr_registers(0)(876) and tmr_registers(1)(876)) or                                            
                            (tmr_registers(1)(876) and tmr_registers(2)(876)) or                                                       
                            (tmr_registers(0)(876) and tmr_registers(2)(876));                                                         
                                                                                                                                     
        global_tmr_voter(1)(877)  <=    (tmr_registers(0)(877) and tmr_registers(1)(877)) or                                            
                            (tmr_registers(1)(877) and tmr_registers(2)(877)) or                                                       
                            (tmr_registers(0)(877) and tmr_registers(2)(877));                                                         
                                                                                                                                     
        global_tmr_voter(1)(878)  <=    (tmr_registers(0)(878) and tmr_registers(1)(878)) or                                            
                            (tmr_registers(1)(878) and tmr_registers(2)(878)) or                                                       
                            (tmr_registers(0)(878) and tmr_registers(2)(878));                                                         
                                                                                                                                     
        global_tmr_voter(1)(879)  <=    (tmr_registers(0)(879) and tmr_registers(1)(879)) or                                            
                            (tmr_registers(1)(879) and tmr_registers(2)(879)) or                                                       
                            (tmr_registers(0)(879) and tmr_registers(2)(879));                                                         
                                                                                                                                     
        global_tmr_voter(1)(880)  <=    (tmr_registers(0)(880) and tmr_registers(1)(880)) or                                            
                            (tmr_registers(1)(880) and tmr_registers(2)(880)) or                                                       
                            (tmr_registers(0)(880) and tmr_registers(2)(880));                                                         
                                                                                                                                     
        global_tmr_voter(1)(881)  <=    (tmr_registers(0)(881) and tmr_registers(1)(881)) or                                            
                            (tmr_registers(1)(881) and tmr_registers(2)(881)) or                                                       
                            (tmr_registers(0)(881) and tmr_registers(2)(881));                                                         
                                                                                                                                     
        global_tmr_voter(1)(882)  <=    (tmr_registers(0)(882) and tmr_registers(1)(882)) or                                            
                            (tmr_registers(1)(882) and tmr_registers(2)(882)) or                                                       
                            (tmr_registers(0)(882) and tmr_registers(2)(882));                                                         
                                                                                                                                     
        global_tmr_voter(1)(883)  <=    (tmr_registers(0)(883) and tmr_registers(1)(883)) or                                            
                            (tmr_registers(1)(883) and tmr_registers(2)(883)) or                                                       
                            (tmr_registers(0)(883) and tmr_registers(2)(883));                                                         
                                                                                                                                     
        global_tmr_voter(1)(884)  <=    (tmr_registers(0)(884) and tmr_registers(1)(884)) or                                            
                            (tmr_registers(1)(884) and tmr_registers(2)(884)) or                                                       
                            (tmr_registers(0)(884) and tmr_registers(2)(884));                                                         
                                                                                                                                     
        global_tmr_voter(1)(885)  <=    (tmr_registers(0)(885) and tmr_registers(1)(885)) or                                            
                            (tmr_registers(1)(885) and tmr_registers(2)(885)) or                                                       
                            (tmr_registers(0)(885) and tmr_registers(2)(885));                                                         
                                                                                                                                     
        global_tmr_voter(1)(886)  <=    (tmr_registers(0)(886) and tmr_registers(1)(886)) or                                            
                            (tmr_registers(1)(886) and tmr_registers(2)(886)) or                                                       
                            (tmr_registers(0)(886) and tmr_registers(2)(886));                                                         
                                                                                                                                     
        global_tmr_voter(1)(887)  <=    (tmr_registers(0)(887) and tmr_registers(1)(887)) or                                            
                            (tmr_registers(1)(887) and tmr_registers(2)(887)) or                                                       
                            (tmr_registers(0)(887) and tmr_registers(2)(887));                                                         
                                                                                                                                     
        global_tmr_voter(1)(888)  <=    (tmr_registers(0)(888) and tmr_registers(1)(888)) or                                            
                            (tmr_registers(1)(888) and tmr_registers(2)(888)) or                                                       
                            (tmr_registers(0)(888) and tmr_registers(2)(888));                                                         
                                                                                                                                     
        global_tmr_voter(1)(889)  <=    (tmr_registers(0)(889) and tmr_registers(1)(889)) or                                            
                            (tmr_registers(1)(889) and tmr_registers(2)(889)) or                                                       
                            (tmr_registers(0)(889) and tmr_registers(2)(889));                                                         
                                                                                                                                     
        global_tmr_voter(1)(890)  <=    (tmr_registers(0)(890) and tmr_registers(1)(890)) or                                            
                            (tmr_registers(1)(890) and tmr_registers(2)(890)) or                                                       
                            (tmr_registers(0)(890) and tmr_registers(2)(890));                                                         
                                                                                                                                     
        global_tmr_voter(1)(891)  <=    (tmr_registers(0)(891) and tmr_registers(1)(891)) or                                            
                            (tmr_registers(1)(891) and tmr_registers(2)(891)) or                                                       
                            (tmr_registers(0)(891) and tmr_registers(2)(891));                                                         
                                                                                                                                     
        global_tmr_voter(1)(892)  <=    (tmr_registers(0)(892) and tmr_registers(1)(892)) or                                            
                            (tmr_registers(1)(892) and tmr_registers(2)(892)) or                                                       
                            (tmr_registers(0)(892) and tmr_registers(2)(892));                                                         
                                                                                                                                     
        global_tmr_voter(1)(893)  <=    (tmr_registers(0)(893) and tmr_registers(1)(893)) or                                            
                            (tmr_registers(1)(893) and tmr_registers(2)(893)) or                                                       
                            (tmr_registers(0)(893) and tmr_registers(2)(893));                                                         
                                                                                                                                     
        global_tmr_voter(1)(894)  <=    (tmr_registers(0)(894) and tmr_registers(1)(894)) or                                            
                            (tmr_registers(1)(894) and tmr_registers(2)(894)) or                                                       
                            (tmr_registers(0)(894) and tmr_registers(2)(894));                                                         
                                                                                                                                     
        global_tmr_voter(1)(895)  <=    (tmr_registers(0)(895) and tmr_registers(1)(895)) or                                            
                            (tmr_registers(1)(895) and tmr_registers(2)(895)) or                                                       
                            (tmr_registers(0)(895) and tmr_registers(2)(895));                                                         
                                                                                                                                     
        global_tmr_voter(1)(896)  <=    (tmr_registers(0)(896) and tmr_registers(1)(896)) or                                            
                            (tmr_registers(1)(896) and tmr_registers(2)(896)) or                                                       
                            (tmr_registers(0)(896) and tmr_registers(2)(896));                                                         
                                                                                                                                     
        global_tmr_voter(1)(897)  <=    (tmr_registers(0)(897) and tmr_registers(1)(897)) or                                            
                            (tmr_registers(1)(897) and tmr_registers(2)(897)) or                                                       
                            (tmr_registers(0)(897) and tmr_registers(2)(897));                                                         
                                                                                                                                     
        global_tmr_voter(1)(898)  <=    (tmr_registers(0)(898) and tmr_registers(1)(898)) or                                            
                            (tmr_registers(1)(898) and tmr_registers(2)(898)) or                                                       
                            (tmr_registers(0)(898) and tmr_registers(2)(898));                                                         
                                                                                                                                     
        global_tmr_voter(1)(899)  <=    (tmr_registers(0)(899) and tmr_registers(1)(899)) or                                            
                            (tmr_registers(1)(899) and tmr_registers(2)(899)) or                                                       
                            (tmr_registers(0)(899) and tmr_registers(2)(899));                                                         
                                                                                                                                     
        global_tmr_voter(1)(900)  <=    (tmr_registers(0)(900) and tmr_registers(1)(900)) or                                            
                            (tmr_registers(1)(900) and tmr_registers(2)(900)) or                                                       
                            (tmr_registers(0)(900) and tmr_registers(2)(900));                                                         
                                                                                                                                     
        global_tmr_voter(1)(901)  <=    (tmr_registers(0)(901) and tmr_registers(1)(901)) or                                            
                            (tmr_registers(1)(901) and tmr_registers(2)(901)) or                                                       
                            (tmr_registers(0)(901) and tmr_registers(2)(901));                                                         
                                                                                                                                     
        global_tmr_voter(1)(902)  <=    (tmr_registers(0)(902) and tmr_registers(1)(902)) or                                            
                            (tmr_registers(1)(902) and tmr_registers(2)(902)) or                                                       
                            (tmr_registers(0)(902) and tmr_registers(2)(902));                                                         
                                                                                                                                     
        global_tmr_voter(1)(903)  <=    (tmr_registers(0)(903) and tmr_registers(1)(903)) or                                            
                            (tmr_registers(1)(903) and tmr_registers(2)(903)) or                                                       
                            (tmr_registers(0)(903) and tmr_registers(2)(903));                                                         
                                                                                                                                     
        global_tmr_voter(1)(904)  <=    (tmr_registers(0)(904) and tmr_registers(1)(904)) or                                            
                            (tmr_registers(1)(904) and tmr_registers(2)(904)) or                                                       
                            (tmr_registers(0)(904) and tmr_registers(2)(904));                                                         
                                                                                                                                     
        global_tmr_voter(1)(905)  <=    (tmr_registers(0)(905) and tmr_registers(1)(905)) or                                            
                            (tmr_registers(1)(905) and tmr_registers(2)(905)) or                                                       
                            (tmr_registers(0)(905) and tmr_registers(2)(905));                                                         
                                                                                                                                     
        global_tmr_voter(1)(906)  <=    (tmr_registers(0)(906) and tmr_registers(1)(906)) or                                            
                            (tmr_registers(1)(906) and tmr_registers(2)(906)) or                                                       
                            (tmr_registers(0)(906) and tmr_registers(2)(906));                                                         
                                                                                                                                     
        global_tmr_voter(1)(907)  <=    (tmr_registers(0)(907) and tmr_registers(1)(907)) or                                            
                            (tmr_registers(1)(907) and tmr_registers(2)(907)) or                                                       
                            (tmr_registers(0)(907) and tmr_registers(2)(907));                                                         
                                                                                                                                     
        global_tmr_voter(1)(908)  <=    (tmr_registers(0)(908) and tmr_registers(1)(908)) or                                            
                            (tmr_registers(1)(908) and tmr_registers(2)(908)) or                                                       
                            (tmr_registers(0)(908) and tmr_registers(2)(908));                                                         
                                                                                                                                     
        global_tmr_voter(1)(909)  <=    (tmr_registers(0)(909) and tmr_registers(1)(909)) or                                            
                            (tmr_registers(1)(909) and tmr_registers(2)(909)) or                                                       
                            (tmr_registers(0)(909) and tmr_registers(2)(909));                                                         
                                                                                                                                     
        global_tmr_voter(1)(910)  <=    (tmr_registers(0)(910) and tmr_registers(1)(910)) or                                            
                            (tmr_registers(1)(910) and tmr_registers(2)(910)) or                                                       
                            (tmr_registers(0)(910) and tmr_registers(2)(910));                                                         
                                                                                                                                     
        global_tmr_voter(1)(911)  <=    (tmr_registers(0)(911) and tmr_registers(1)(911)) or                                            
                            (tmr_registers(1)(911) and tmr_registers(2)(911)) or                                                       
                            (tmr_registers(0)(911) and tmr_registers(2)(911));                                                         
                                                                                                                                     
        global_tmr_voter(1)(912)  <=    (tmr_registers(0)(912) and tmr_registers(1)(912)) or                                            
                            (tmr_registers(1)(912) and tmr_registers(2)(912)) or                                                       
                            (tmr_registers(0)(912) and tmr_registers(2)(912));                                                         
                                                                                                                                     
        global_tmr_voter(1)(913)  <=    (tmr_registers(0)(913) and tmr_registers(1)(913)) or                                            
                            (tmr_registers(1)(913) and tmr_registers(2)(913)) or                                                       
                            (tmr_registers(0)(913) and tmr_registers(2)(913));                                                         
                                                                                                                                     
        global_tmr_voter(1)(914)  <=    (tmr_registers(0)(914) and tmr_registers(1)(914)) or                                            
                            (tmr_registers(1)(914) and tmr_registers(2)(914)) or                                                       
                            (tmr_registers(0)(914) and tmr_registers(2)(914));                                                         
                                                                                                                                     
        global_tmr_voter(1)(915)  <=    (tmr_registers(0)(915) and tmr_registers(1)(915)) or                                            
                            (tmr_registers(1)(915) and tmr_registers(2)(915)) or                                                       
                            (tmr_registers(0)(915) and tmr_registers(2)(915));                                                         
                                                                                                                                     
        global_tmr_voter(1)(916)  <=    (tmr_registers(0)(916) and tmr_registers(1)(916)) or                                            
                            (tmr_registers(1)(916) and tmr_registers(2)(916)) or                                                       
                            (tmr_registers(0)(916) and tmr_registers(2)(916));                                                         
                                                                                                                                     
        global_tmr_voter(1)(917)  <=    (tmr_registers(0)(917) and tmr_registers(1)(917)) or                                            
                            (tmr_registers(1)(917) and tmr_registers(2)(917)) or                                                       
                            (tmr_registers(0)(917) and tmr_registers(2)(917));                                                         
                                                                                                                                     
        global_tmr_voter(1)(918)  <=    (tmr_registers(0)(918) and tmr_registers(1)(918)) or                                            
                            (tmr_registers(1)(918) and tmr_registers(2)(918)) or                                                       
                            (tmr_registers(0)(918) and tmr_registers(2)(918));                                                         
                                                                                                                                     
        global_tmr_voter(1)(919)  <=    (tmr_registers(0)(919) and tmr_registers(1)(919)) or                                            
                            (tmr_registers(1)(919) and tmr_registers(2)(919)) or                                                       
                            (tmr_registers(0)(919) and tmr_registers(2)(919));                                                         
                                                                                                                                     
        global_tmr_voter(1)(920)  <=    (tmr_registers(0)(920) and tmr_registers(1)(920)) or                                            
                            (tmr_registers(1)(920) and tmr_registers(2)(920)) or                                                       
                            (tmr_registers(0)(920) and tmr_registers(2)(920));                                                         
                                                                                                                                     
        global_tmr_voter(1)(921)  <=    (tmr_registers(0)(921) and tmr_registers(1)(921)) or                                            
                            (tmr_registers(1)(921) and tmr_registers(2)(921)) or                                                       
                            (tmr_registers(0)(921) and tmr_registers(2)(921));                                                         
                                                                                                                                     
        global_tmr_voter(1)(922)  <=    (tmr_registers(0)(922) and tmr_registers(1)(922)) or                                            
                            (tmr_registers(1)(922) and tmr_registers(2)(922)) or                                                       
                            (tmr_registers(0)(922) and tmr_registers(2)(922));                                                         
                                                                                                                                     
        global_tmr_voter(1)(923)  <=    (tmr_registers(0)(923) and tmr_registers(1)(923)) or                                            
                            (tmr_registers(1)(923) and tmr_registers(2)(923)) or                                                       
                            (tmr_registers(0)(923) and tmr_registers(2)(923));                                                         
                                                                                                                                     
        global_tmr_voter(1)(924)  <=    (tmr_registers(0)(924) and tmr_registers(1)(924)) or                                            
                            (tmr_registers(1)(924) and tmr_registers(2)(924)) or                                                       
                            (tmr_registers(0)(924) and tmr_registers(2)(924));                                                         
                                                                                                                                     
        global_tmr_voter(1)(925)  <=    (tmr_registers(0)(925) and tmr_registers(1)(925)) or                                            
                            (tmr_registers(1)(925) and tmr_registers(2)(925)) or                                                       
                            (tmr_registers(0)(925) and tmr_registers(2)(925));                                                         
                                                                                                                                     
        global_tmr_voter(1)(926)  <=    (tmr_registers(0)(926) and tmr_registers(1)(926)) or                                            
                            (tmr_registers(1)(926) and tmr_registers(2)(926)) or                                                       
                            (tmr_registers(0)(926) and tmr_registers(2)(926));                                                         
                                                                                                                                     
        global_tmr_voter(1)(927)  <=    (tmr_registers(0)(927) and tmr_registers(1)(927)) or                                            
                            (tmr_registers(1)(927) and tmr_registers(2)(927)) or                                                       
                            (tmr_registers(0)(927) and tmr_registers(2)(927));                                                         
                                                                                                                                     
        global_tmr_voter(1)(928)  <=    (tmr_registers(0)(928) and tmr_registers(1)(928)) or                                            
                            (tmr_registers(1)(928) and tmr_registers(2)(928)) or                                                       
                            (tmr_registers(0)(928) and tmr_registers(2)(928));                                                         
                                                                                                                                     
        global_tmr_voter(1)(929)  <=    (tmr_registers(0)(929) and tmr_registers(1)(929)) or                                            
                            (tmr_registers(1)(929) and tmr_registers(2)(929)) or                                                       
                            (tmr_registers(0)(929) and tmr_registers(2)(929));                                                         
                                                                                                                                     
        global_tmr_voter(1)(930)  <=    (tmr_registers(0)(930) and tmr_registers(1)(930)) or                                            
                            (tmr_registers(1)(930) and tmr_registers(2)(930)) or                                                       
                            (tmr_registers(0)(930) and tmr_registers(2)(930));                                                         
                                                                                                                                     
        global_tmr_voter(1)(931)  <=    (tmr_registers(0)(931) and tmr_registers(1)(931)) or                                            
                            (tmr_registers(1)(931) and tmr_registers(2)(931)) or                                                       
                            (tmr_registers(0)(931) and tmr_registers(2)(931));                                                         
                                                                                                                                     
        global_tmr_voter(1)(932)  <=    (tmr_registers(0)(932) and tmr_registers(1)(932)) or                                            
                            (tmr_registers(1)(932) and tmr_registers(2)(932)) or                                                       
                            (tmr_registers(0)(932) and tmr_registers(2)(932));                                                         
                                                                                                                                     
        global_tmr_voter(1)(933)  <=    (tmr_registers(0)(933) and tmr_registers(1)(933)) or                                            
                            (tmr_registers(1)(933) and tmr_registers(2)(933)) or                                                       
                            (tmr_registers(0)(933) and tmr_registers(2)(933));                                                         
                                                                                                                                     
        global_tmr_voter(1)(934)  <=    (tmr_registers(0)(934) and tmr_registers(1)(934)) or                                            
                            (tmr_registers(1)(934) and tmr_registers(2)(934)) or                                                       
                            (tmr_registers(0)(934) and tmr_registers(2)(934));                                                         
                                                                                                                                     
        global_tmr_voter(1)(935)  <=    (tmr_registers(0)(935) and tmr_registers(1)(935)) or                                            
                            (tmr_registers(1)(935) and tmr_registers(2)(935)) or                                                       
                            (tmr_registers(0)(935) and tmr_registers(2)(935));                                                         
                                                                                                                                     
        global_tmr_voter(1)(936)  <=    (tmr_registers(0)(936) and tmr_registers(1)(936)) or                                            
                            (tmr_registers(1)(936) and tmr_registers(2)(936)) or                                                       
                            (tmr_registers(0)(936) and tmr_registers(2)(936));                                                         
                                                                                                                                     
        global_tmr_voter(1)(937)  <=    (tmr_registers(0)(937) and tmr_registers(1)(937)) or                                            
                            (tmr_registers(1)(937) and tmr_registers(2)(937)) or                                                       
                            (tmr_registers(0)(937) and tmr_registers(2)(937));                                                         
                                                                                                                                     
        global_tmr_voter(1)(938)  <=    (tmr_registers(0)(938) and tmr_registers(1)(938)) or                                            
                            (tmr_registers(1)(938) and tmr_registers(2)(938)) or                                                       
                            (tmr_registers(0)(938) and tmr_registers(2)(938));                                                         
                                                                                                                                     
        global_tmr_voter(1)(939)  <=    (tmr_registers(0)(939) and tmr_registers(1)(939)) or                                            
                            (tmr_registers(1)(939) and tmr_registers(2)(939)) or                                                       
                            (tmr_registers(0)(939) and tmr_registers(2)(939));                                                         
                                                                                                                                     
        global_tmr_voter(1)(940)  <=    (tmr_registers(0)(940) and tmr_registers(1)(940)) or                                            
                            (tmr_registers(1)(940) and tmr_registers(2)(940)) or                                                       
                            (tmr_registers(0)(940) and tmr_registers(2)(940));                                                         
                                                                                                                                     
        global_tmr_voter(1)(941)  <=    (tmr_registers(0)(941) and tmr_registers(1)(941)) or                                            
                            (tmr_registers(1)(941) and tmr_registers(2)(941)) or                                                       
                            (tmr_registers(0)(941) and tmr_registers(2)(941));                                                         
                                                                                                                                     
        global_tmr_voter(1)(942)  <=    (tmr_registers(0)(942) and tmr_registers(1)(942)) or                                            
                            (tmr_registers(1)(942) and tmr_registers(2)(942)) or                                                       
                            (tmr_registers(0)(942) and tmr_registers(2)(942));                                                         
                                                                                                                                     
        global_tmr_voter(1)(943)  <=    (tmr_registers(0)(943) and tmr_registers(1)(943)) or                                            
                            (tmr_registers(1)(943) and tmr_registers(2)(943)) or                                                       
                            (tmr_registers(0)(943) and tmr_registers(2)(943));                                                         
                                                                                                                                     
        global_tmr_voter(1)(944)  <=    (tmr_registers(0)(944) and tmr_registers(1)(944)) or                                            
                            (tmr_registers(1)(944) and tmr_registers(2)(944)) or                                                       
                            (tmr_registers(0)(944) and tmr_registers(2)(944));                                                         
                                                                                                                                     
        global_tmr_voter(1)(945)  <=    (tmr_registers(0)(945) and tmr_registers(1)(945)) or                                            
                            (tmr_registers(1)(945) and tmr_registers(2)(945)) or                                                       
                            (tmr_registers(0)(945) and tmr_registers(2)(945));                                                         
                                                                                                                                     
        global_tmr_voter(1)(946)  <=    (tmr_registers(0)(946) and tmr_registers(1)(946)) or                                            
                            (tmr_registers(1)(946) and tmr_registers(2)(946)) or                                                       
                            (tmr_registers(0)(946) and tmr_registers(2)(946));                                                         
                                                                                                                                     
        global_tmr_voter(1)(947)  <=    (tmr_registers(0)(947) and tmr_registers(1)(947)) or                                            
                            (tmr_registers(1)(947) and tmr_registers(2)(947)) or                                                       
                            (tmr_registers(0)(947) and tmr_registers(2)(947));                                                         
                                                                                                                                     
        global_tmr_voter(1)(948)  <=    (tmr_registers(0)(948) and tmr_registers(1)(948)) or                                            
                            (tmr_registers(1)(948) and tmr_registers(2)(948)) or                                                       
                            (tmr_registers(0)(948) and tmr_registers(2)(948));                                                         
                                                                                                                                     
        global_tmr_voter(1)(949)  <=    (tmr_registers(0)(949) and tmr_registers(1)(949)) or                                            
                            (tmr_registers(1)(949) and tmr_registers(2)(949)) or                                                       
                            (tmr_registers(0)(949) and tmr_registers(2)(949));                                                         
                                                                                                                                     
        global_tmr_voter(1)(950)  <=    (tmr_registers(0)(950) and tmr_registers(1)(950)) or                                            
                            (tmr_registers(1)(950) and tmr_registers(2)(950)) or                                                       
                            (tmr_registers(0)(950) and tmr_registers(2)(950));                                                         
                                                                                                                                     
        global_tmr_voter(1)(951)  <=    (tmr_registers(0)(951) and tmr_registers(1)(951)) or                                            
                            (tmr_registers(1)(951) and tmr_registers(2)(951)) or                                                       
                            (tmr_registers(0)(951) and tmr_registers(2)(951));                                                         
                                                                                                                                     
        global_tmr_voter(1)(952)  <=    (tmr_registers(0)(952) and tmr_registers(1)(952)) or                                            
                            (tmr_registers(1)(952) and tmr_registers(2)(952)) or                                                       
                            (tmr_registers(0)(952) and tmr_registers(2)(952));                                                         
                                                                                                                                     
        global_tmr_voter(1)(953)  <=    (tmr_registers(0)(953) and tmr_registers(1)(953)) or                                            
                            (tmr_registers(1)(953) and tmr_registers(2)(953)) or                                                       
                            (tmr_registers(0)(953) and tmr_registers(2)(953));                                                         
                                                                                                                                     
        global_tmr_voter(1)(954)  <=    (tmr_registers(0)(954) and tmr_registers(1)(954)) or                                            
                            (tmr_registers(1)(954) and tmr_registers(2)(954)) or                                                       
                            (tmr_registers(0)(954) and tmr_registers(2)(954));                                                         
                                                                                                                                     
        global_tmr_voter(1)(955)  <=    (tmr_registers(0)(955) and tmr_registers(1)(955)) or                                            
                            (tmr_registers(1)(955) and tmr_registers(2)(955)) or                                                       
                            (tmr_registers(0)(955) and tmr_registers(2)(955));                                                         
                                                                                                                                     
        global_tmr_voter(1)(956)  <=    (tmr_registers(0)(956) and tmr_registers(1)(956)) or                                            
                            (tmr_registers(1)(956) and tmr_registers(2)(956)) or                                                       
                            (tmr_registers(0)(956) and tmr_registers(2)(956));                                                         
                                                                                                                                     
        global_tmr_voter(1)(957)  <=    (tmr_registers(0)(957) and tmr_registers(1)(957)) or                                            
                            (tmr_registers(1)(957) and tmr_registers(2)(957)) or                                                       
                            (tmr_registers(0)(957) and tmr_registers(2)(957));                                                         
                                                                                                                                     
        global_tmr_voter(1)(958)  <=    (tmr_registers(0)(958) and tmr_registers(1)(958)) or                                            
                            (tmr_registers(1)(958) and tmr_registers(2)(958)) or                                                       
                            (tmr_registers(0)(958) and tmr_registers(2)(958));                                                         
                                                                                                                                     
        global_tmr_voter(1)(959)  <=    (tmr_registers(0)(959) and tmr_registers(1)(959)) or                                            
                            (tmr_registers(1)(959) and tmr_registers(2)(959)) or                                                       
                            (tmr_registers(0)(959) and tmr_registers(2)(959));                                                         
                                                                                                                                     
        global_tmr_voter(1)(960)  <=    (tmr_registers(0)(960) and tmr_registers(1)(960)) or                                            
                            (tmr_registers(1)(960) and tmr_registers(2)(960)) or                                                       
                            (tmr_registers(0)(960) and tmr_registers(2)(960));                                                         
                                                                                                                                     
        global_tmr_voter(1)(961)  <=    (tmr_registers(0)(961) and tmr_registers(1)(961)) or                                            
                            (tmr_registers(1)(961) and tmr_registers(2)(961)) or                                                       
                            (tmr_registers(0)(961) and tmr_registers(2)(961));                                                         
                                                                                                                                     
        global_tmr_voter(1)(962)  <=    (tmr_registers(0)(962) and tmr_registers(1)(962)) or                                            
                            (tmr_registers(1)(962) and tmr_registers(2)(962)) or                                                       
                            (tmr_registers(0)(962) and tmr_registers(2)(962));                                                         
                                                                                                                                     
        global_tmr_voter(1)(963)  <=    (tmr_registers(0)(963) and tmr_registers(1)(963)) or                                            
                            (tmr_registers(1)(963) and tmr_registers(2)(963)) or                                                       
                            (tmr_registers(0)(963) and tmr_registers(2)(963));                                                         
                                                                                                                                     
        global_tmr_voter(1)(964)  <=    (tmr_registers(0)(964) and tmr_registers(1)(964)) or                                            
                            (tmr_registers(1)(964) and tmr_registers(2)(964)) or                                                       
                            (tmr_registers(0)(964) and tmr_registers(2)(964));                                                         
                                                                                                                                     
        global_tmr_voter(1)(965)  <=    (tmr_registers(0)(965) and tmr_registers(1)(965)) or                                            
                            (tmr_registers(1)(965) and tmr_registers(2)(965)) or                                                       
                            (tmr_registers(0)(965) and tmr_registers(2)(965));                                                         
                                                                                                                                     
        global_tmr_voter(1)(966)  <=    (tmr_registers(0)(966) and tmr_registers(1)(966)) or                                            
                            (tmr_registers(1)(966) and tmr_registers(2)(966)) or                                                       
                            (tmr_registers(0)(966) and tmr_registers(2)(966));                                                         
                                                                                                                                     
        global_tmr_voter(1)(967)  <=    (tmr_registers(0)(967) and tmr_registers(1)(967)) or                                            
                            (tmr_registers(1)(967) and tmr_registers(2)(967)) or                                                       
                            (tmr_registers(0)(967) and tmr_registers(2)(967));                                                         
                                                                                                                                     
        global_tmr_voter(1)(968)  <=    (tmr_registers(0)(968) and tmr_registers(1)(968)) or                                            
                            (tmr_registers(1)(968) and tmr_registers(2)(968)) or                                                       
                            (tmr_registers(0)(968) and tmr_registers(2)(968));                                                         
                                                                                                                                     
        global_tmr_voter(1)(969)  <=    (tmr_registers(0)(969) and tmr_registers(1)(969)) or                                            
                            (tmr_registers(1)(969) and tmr_registers(2)(969)) or                                                       
                            (tmr_registers(0)(969) and tmr_registers(2)(969));                                                         
                                                                                                                                     
        global_tmr_voter(1)(970)  <=    (tmr_registers(0)(970) and tmr_registers(1)(970)) or                                            
                            (tmr_registers(1)(970) and tmr_registers(2)(970)) or                                                       
                            (tmr_registers(0)(970) and tmr_registers(2)(970));                                                         
                                                                                                                                     
        global_tmr_voter(1)(971)  <=    (tmr_registers(0)(971) and tmr_registers(1)(971)) or                                            
                            (tmr_registers(1)(971) and tmr_registers(2)(971)) or                                                       
                            (tmr_registers(0)(971) and tmr_registers(2)(971));                                                         
                                                                                                                                     
        global_tmr_voter(1)(972)  <=    (tmr_registers(0)(972) and tmr_registers(1)(972)) or                                            
                            (tmr_registers(1)(972) and tmr_registers(2)(972)) or                                                       
                            (tmr_registers(0)(972) and tmr_registers(2)(972));                                                         
                                                                                                                                     
        global_tmr_voter(1)(973)  <=    (tmr_registers(0)(973) and tmr_registers(1)(973)) or                                            
                            (tmr_registers(1)(973) and tmr_registers(2)(973)) or                                                       
                            (tmr_registers(0)(973) and tmr_registers(2)(973));                                                         
                                                                                                                                     
        global_tmr_voter(1)(974)  <=    (tmr_registers(0)(974) and tmr_registers(1)(974)) or                                            
                            (tmr_registers(1)(974) and tmr_registers(2)(974)) or                                                       
                            (tmr_registers(0)(974) and tmr_registers(2)(974));                                                         
                                                                                                                                     
        global_tmr_voter(1)(975)  <=    (tmr_registers(0)(975) and tmr_registers(1)(975)) or                                            
                            (tmr_registers(1)(975) and tmr_registers(2)(975)) or                                                       
                            (tmr_registers(0)(975) and tmr_registers(2)(975));                                                         
                                                                                                                                     
        global_tmr_voter(1)(976)  <=    (tmr_registers(0)(976) and tmr_registers(1)(976)) or                                            
                            (tmr_registers(1)(976) and tmr_registers(2)(976)) or                                                       
                            (tmr_registers(0)(976) and tmr_registers(2)(976));                                                         
                                                                                                                                     
        global_tmr_voter(1)(977)  <=    (tmr_registers(0)(977) and tmr_registers(1)(977)) or                                            
                            (tmr_registers(1)(977) and tmr_registers(2)(977)) or                                                       
                            (tmr_registers(0)(977) and tmr_registers(2)(977));                                                         
                                                                                                                                     
        global_tmr_voter(1)(978)  <=    (tmr_registers(0)(978) and tmr_registers(1)(978)) or                                            
                            (tmr_registers(1)(978) and tmr_registers(2)(978)) or                                                       
                            (tmr_registers(0)(978) and tmr_registers(2)(978));                                                         
                                                                                                                                     
        global_tmr_voter(1)(979)  <=    (tmr_registers(0)(979) and tmr_registers(1)(979)) or                                            
                            (tmr_registers(1)(979) and tmr_registers(2)(979)) or                                                       
                            (tmr_registers(0)(979) and tmr_registers(2)(979));                                                         
                                                                                                                                     
        global_tmr_voter(1)(980)  <=    (tmr_registers(0)(980) and tmr_registers(1)(980)) or                                            
                            (tmr_registers(1)(980) and tmr_registers(2)(980)) or                                                       
                            (tmr_registers(0)(980) and tmr_registers(2)(980));                                                         
                                                                                                                                     
        global_tmr_voter(1)(981)  <=    (tmr_registers(0)(981) and tmr_registers(1)(981)) or                                            
                            (tmr_registers(1)(981) and tmr_registers(2)(981)) or                                                       
                            (tmr_registers(0)(981) and tmr_registers(2)(981));                                                         
                                                                                                                                     
        global_tmr_voter(1)(982)  <=    (tmr_registers(0)(982) and tmr_registers(1)(982)) or                                            
                            (tmr_registers(1)(982) and tmr_registers(2)(982)) or                                                       
                            (tmr_registers(0)(982) and tmr_registers(2)(982));                                                         
                                                                                                                                     
        global_tmr_voter(1)(983)  <=    (tmr_registers(0)(983) and tmr_registers(1)(983)) or                                            
                            (tmr_registers(1)(983) and tmr_registers(2)(983)) or                                                       
                            (tmr_registers(0)(983) and tmr_registers(2)(983));                                                         
                                                                                                                                     
        global_tmr_voter(1)(984)  <=    (tmr_registers(0)(984) and tmr_registers(1)(984)) or                                            
                            (tmr_registers(1)(984) and tmr_registers(2)(984)) or                                                       
                            (tmr_registers(0)(984) and tmr_registers(2)(984));                                                         
                                                                                                                                     
        global_tmr_voter(1)(985)  <=    (tmr_registers(0)(985) and tmr_registers(1)(985)) or                                            
                            (tmr_registers(1)(985) and tmr_registers(2)(985)) or                                                       
                            (tmr_registers(0)(985) and tmr_registers(2)(985));                                                         
                                                                                                                                     
        global_tmr_voter(1)(986)  <=    (tmr_registers(0)(986) and tmr_registers(1)(986)) or                                            
                            (tmr_registers(1)(986) and tmr_registers(2)(986)) or                                                       
                            (tmr_registers(0)(986) and tmr_registers(2)(986));                                                         
                                                                                                                                     
        global_tmr_voter(1)(987)  <=    (tmr_registers(0)(987) and tmr_registers(1)(987)) or                                            
                            (tmr_registers(1)(987) and tmr_registers(2)(987)) or                                                       
                            (tmr_registers(0)(987) and tmr_registers(2)(987));                                                         
                                                                                                                                     
        global_tmr_voter(1)(988)  <=    (tmr_registers(0)(988) and tmr_registers(1)(988)) or                                            
                            (tmr_registers(1)(988) and tmr_registers(2)(988)) or                                                       
                            (tmr_registers(0)(988) and tmr_registers(2)(988));                                                         
                                                                                                                                     
        global_tmr_voter(1)(989)  <=    (tmr_registers(0)(989) and tmr_registers(1)(989)) or                                            
                            (tmr_registers(1)(989) and tmr_registers(2)(989)) or                                                       
                            (tmr_registers(0)(989) and tmr_registers(2)(989));                                                         
                                                                                                                                     
        global_tmr_voter(1)(990)  <=    (tmr_registers(0)(990) and tmr_registers(1)(990)) or                                            
                            (tmr_registers(1)(990) and tmr_registers(2)(990)) or                                                       
                            (tmr_registers(0)(990) and tmr_registers(2)(990));                                                         
                                                                                                                                     
        global_tmr_voter(1)(991)  <=    (tmr_registers(0)(991) and tmr_registers(1)(991)) or                                            
                            (tmr_registers(1)(991) and tmr_registers(2)(991)) or                                                       
                            (tmr_registers(0)(991) and tmr_registers(2)(991));                                                         
                                                                                                                                     
        global_tmr_voter(1)(992)  <=    (tmr_registers(0)(992) and tmr_registers(1)(992)) or                                            
                            (tmr_registers(1)(992) and tmr_registers(2)(992)) or                                                       
                            (tmr_registers(0)(992) and tmr_registers(2)(992));                                                         
                                                                                                                                     
        global_tmr_voter(1)(993)  <=    (tmr_registers(0)(993) and tmr_registers(1)(993)) or                                            
                            (tmr_registers(1)(993) and tmr_registers(2)(993)) or                                                       
                            (tmr_registers(0)(993) and tmr_registers(2)(993));                                                         
                                                                                                                                     
        global_tmr_voter(1)(994)  <=    (tmr_registers(0)(994) and tmr_registers(1)(994)) or                                            
                            (tmr_registers(1)(994) and tmr_registers(2)(994)) or                                                       
                            (tmr_registers(0)(994) and tmr_registers(2)(994));                                                         
                                                                                                                                     
        global_tmr_voter(1)(995)  <=    (tmr_registers(0)(995) and tmr_registers(1)(995)) or                                            
                            (tmr_registers(1)(995) and tmr_registers(2)(995)) or                                                       
                            (tmr_registers(0)(995) and tmr_registers(2)(995));                                                         
                                                                                                                                     
        global_tmr_voter(1)(996)  <=    (tmr_registers(0)(996) and tmr_registers(1)(996)) or                                            
                            (tmr_registers(1)(996) and tmr_registers(2)(996)) or                                                       
                            (tmr_registers(0)(996) and tmr_registers(2)(996));                                                         
                                                                                                                                     
        global_tmr_voter(1)(997)  <=    (tmr_registers(0)(997) and tmr_registers(1)(997)) or                                            
                            (tmr_registers(1)(997) and tmr_registers(2)(997)) or                                                       
                            (tmr_registers(0)(997) and tmr_registers(2)(997));                                                         
                                                                                                                                     
        global_tmr_voter(1)(998)  <=    (tmr_registers(0)(998) and tmr_registers(1)(998)) or                                            
                            (tmr_registers(1)(998) and tmr_registers(2)(998)) or                                                       
                            (tmr_registers(0)(998) and tmr_registers(2)(998));                                                         
                                                                                                                                     
        global_tmr_voter(1)(999)  <=    (tmr_registers(0)(999) and tmr_registers(1)(999)) or                                            
                            (tmr_registers(1)(999) and tmr_registers(2)(999)) or                                                       
                            (tmr_registers(0)(999) and tmr_registers(2)(999));                                                         
                                                                                                                                     
        global_tmr_voter(2)(1)  <=    (tmr_registers(0)(1) and tmr_registers(1)(1)) or                                            
                            (tmr_registers(1)(1) and tmr_registers(2)(1)) or                                                       
                            (tmr_registers(0)(1) and tmr_registers(2)(1));                                                         
                                                                                                                                     
        global_tmr_voter(2)(2)  <=    (tmr_registers(0)(2) and tmr_registers(1)(2)) or                                            
                            (tmr_registers(1)(2) and tmr_registers(2)(2)) or                                                       
                            (tmr_registers(0)(2) and tmr_registers(2)(2));                                                         
                                                                                                                                     
        global_tmr_voter(2)(3)  <=    (tmr_registers(0)(3) and tmr_registers(1)(3)) or                                            
                            (tmr_registers(1)(3) and tmr_registers(2)(3)) or                                                       
                            (tmr_registers(0)(3) and tmr_registers(2)(3));                                                         
                                                                                                                                     
        global_tmr_voter(2)(4)  <=    (tmr_registers(0)(4) and tmr_registers(1)(4)) or                                            
                            (tmr_registers(1)(4) and tmr_registers(2)(4)) or                                                       
                            (tmr_registers(0)(4) and tmr_registers(2)(4));                                                         
                                                                                                                                     
        global_tmr_voter(2)(5)  <=    (tmr_registers(0)(5) and tmr_registers(1)(5)) or                                            
                            (tmr_registers(1)(5) and tmr_registers(2)(5)) or                                                       
                            (tmr_registers(0)(5) and tmr_registers(2)(5));                                                         
                                                                                                                                     
        global_tmr_voter(2)(6)  <=    (tmr_registers(0)(6) and tmr_registers(1)(6)) or                                            
                            (tmr_registers(1)(6) and tmr_registers(2)(6)) or                                                       
                            (tmr_registers(0)(6) and tmr_registers(2)(6));                                                         
                                                                                                                                     
        global_tmr_voter(2)(7)  <=    (tmr_registers(0)(7) and tmr_registers(1)(7)) or                                            
                            (tmr_registers(1)(7) and tmr_registers(2)(7)) or                                                       
                            (tmr_registers(0)(7) and tmr_registers(2)(7));                                                         
                                                                                                                                     
        global_tmr_voter(2)(8)  <=    (tmr_registers(0)(8) and tmr_registers(1)(8)) or                                            
                            (tmr_registers(1)(8) and tmr_registers(2)(8)) or                                                       
                            (tmr_registers(0)(8) and tmr_registers(2)(8));                                                         
                                                                                                                                     
        global_tmr_voter(2)(9)  <=    (tmr_registers(0)(9) and tmr_registers(1)(9)) or                                            
                            (tmr_registers(1)(9) and tmr_registers(2)(9)) or                                                       
                            (tmr_registers(0)(9) and tmr_registers(2)(9));                                                         
                                                                                                                                     
        global_tmr_voter(2)(10)  <=    (tmr_registers(0)(10) and tmr_registers(1)(10)) or                                            
                            (tmr_registers(1)(10) and tmr_registers(2)(10)) or                                                       
                            (tmr_registers(0)(10) and tmr_registers(2)(10));                                                         
                                                                                                                                     
        global_tmr_voter(2)(11)  <=    (tmr_registers(0)(11) and tmr_registers(1)(11)) or                                            
                            (tmr_registers(1)(11) and tmr_registers(2)(11)) or                                                       
                            (tmr_registers(0)(11) and tmr_registers(2)(11));                                                         
                                                                                                                                     
        global_tmr_voter(2)(12)  <=    (tmr_registers(0)(12) and tmr_registers(1)(12)) or                                            
                            (tmr_registers(1)(12) and tmr_registers(2)(12)) or                                                       
                            (tmr_registers(0)(12) and tmr_registers(2)(12));                                                         
                                                                                                                                     
        global_tmr_voter(2)(13)  <=    (tmr_registers(0)(13) and tmr_registers(1)(13)) or                                            
                            (tmr_registers(1)(13) and tmr_registers(2)(13)) or                                                       
                            (tmr_registers(0)(13) and tmr_registers(2)(13));                                                         
                                                                                                                                     
        global_tmr_voter(2)(14)  <=    (tmr_registers(0)(14) and tmr_registers(1)(14)) or                                            
                            (tmr_registers(1)(14) and tmr_registers(2)(14)) or                                                       
                            (tmr_registers(0)(14) and tmr_registers(2)(14));                                                         
                                                                                                                                     
        global_tmr_voter(2)(15)  <=    (tmr_registers(0)(15) and tmr_registers(1)(15)) or                                            
                            (tmr_registers(1)(15) and tmr_registers(2)(15)) or                                                       
                            (tmr_registers(0)(15) and tmr_registers(2)(15));                                                         
                                                                                                                                     
        global_tmr_voter(2)(16)  <=    (tmr_registers(0)(16) and tmr_registers(1)(16)) or                                            
                            (tmr_registers(1)(16) and tmr_registers(2)(16)) or                                                       
                            (tmr_registers(0)(16) and tmr_registers(2)(16));                                                         
                                                                                                                                     
        global_tmr_voter(2)(17)  <=    (tmr_registers(0)(17) and tmr_registers(1)(17)) or                                            
                            (tmr_registers(1)(17) and tmr_registers(2)(17)) or                                                       
                            (tmr_registers(0)(17) and tmr_registers(2)(17));                                                         
                                                                                                                                     
        global_tmr_voter(2)(18)  <=    (tmr_registers(0)(18) and tmr_registers(1)(18)) or                                            
                            (tmr_registers(1)(18) and tmr_registers(2)(18)) or                                                       
                            (tmr_registers(0)(18) and tmr_registers(2)(18));                                                         
                                                                                                                                     
        global_tmr_voter(2)(19)  <=    (tmr_registers(0)(19) and tmr_registers(1)(19)) or                                            
                            (tmr_registers(1)(19) and tmr_registers(2)(19)) or                                                       
                            (tmr_registers(0)(19) and tmr_registers(2)(19));                                                         
                                                                                                                                     
        global_tmr_voter(2)(20)  <=    (tmr_registers(0)(20) and tmr_registers(1)(20)) or                                            
                            (tmr_registers(1)(20) and tmr_registers(2)(20)) or                                                       
                            (tmr_registers(0)(20) and tmr_registers(2)(20));                                                         
                                                                                                                                     
        global_tmr_voter(2)(21)  <=    (tmr_registers(0)(21) and tmr_registers(1)(21)) or                                            
                            (tmr_registers(1)(21) and tmr_registers(2)(21)) or                                                       
                            (tmr_registers(0)(21) and tmr_registers(2)(21));                                                         
                                                                                                                                     
        global_tmr_voter(2)(22)  <=    (tmr_registers(0)(22) and tmr_registers(1)(22)) or                                            
                            (tmr_registers(1)(22) and tmr_registers(2)(22)) or                                                       
                            (tmr_registers(0)(22) and tmr_registers(2)(22));                                                         
                                                                                                                                     
        global_tmr_voter(2)(23)  <=    (tmr_registers(0)(23) and tmr_registers(1)(23)) or                                            
                            (tmr_registers(1)(23) and tmr_registers(2)(23)) or                                                       
                            (tmr_registers(0)(23) and tmr_registers(2)(23));                                                         
                                                                                                                                     
        global_tmr_voter(2)(24)  <=    (tmr_registers(0)(24) and tmr_registers(1)(24)) or                                            
                            (tmr_registers(1)(24) and tmr_registers(2)(24)) or                                                       
                            (tmr_registers(0)(24) and tmr_registers(2)(24));                                                         
                                                                                                                                     
        global_tmr_voter(2)(25)  <=    (tmr_registers(0)(25) and tmr_registers(1)(25)) or                                            
                            (tmr_registers(1)(25) and tmr_registers(2)(25)) or                                                       
                            (tmr_registers(0)(25) and tmr_registers(2)(25));                                                         
                                                                                                                                     
        global_tmr_voter(2)(26)  <=    (tmr_registers(0)(26) and tmr_registers(1)(26)) or                                            
                            (tmr_registers(1)(26) and tmr_registers(2)(26)) or                                                       
                            (tmr_registers(0)(26) and tmr_registers(2)(26));                                                         
                                                                                                                                     
        global_tmr_voter(2)(27)  <=    (tmr_registers(0)(27) and tmr_registers(1)(27)) or                                            
                            (tmr_registers(1)(27) and tmr_registers(2)(27)) or                                                       
                            (tmr_registers(0)(27) and tmr_registers(2)(27));                                                         
                                                                                                                                     
        global_tmr_voter(2)(28)  <=    (tmr_registers(0)(28) and tmr_registers(1)(28)) or                                            
                            (tmr_registers(1)(28) and tmr_registers(2)(28)) or                                                       
                            (tmr_registers(0)(28) and tmr_registers(2)(28));                                                         
                                                                                                                                     
        global_tmr_voter(2)(29)  <=    (tmr_registers(0)(29) and tmr_registers(1)(29)) or                                            
                            (tmr_registers(1)(29) and tmr_registers(2)(29)) or                                                       
                            (tmr_registers(0)(29) and tmr_registers(2)(29));                                                         
                                                                                                                                     
        global_tmr_voter(2)(30)  <=    (tmr_registers(0)(30) and tmr_registers(1)(30)) or                                            
                            (tmr_registers(1)(30) and tmr_registers(2)(30)) or                                                       
                            (tmr_registers(0)(30) and tmr_registers(2)(30));                                                         
                                                                                                                                     
        global_tmr_voter(2)(31)  <=    (tmr_registers(0)(31) and tmr_registers(1)(31)) or                                            
                            (tmr_registers(1)(31) and tmr_registers(2)(31)) or                                                       
                            (tmr_registers(0)(31) and tmr_registers(2)(31));                                                         
                                                                                                                                     
        global_tmr_voter(2)(32)  <=    (tmr_registers(0)(32) and tmr_registers(1)(32)) or                                            
                            (tmr_registers(1)(32) and tmr_registers(2)(32)) or                                                       
                            (tmr_registers(0)(32) and tmr_registers(2)(32));                                                         
                                                                                                                                     
        global_tmr_voter(2)(33)  <=    (tmr_registers(0)(33) and tmr_registers(1)(33)) or                                            
                            (tmr_registers(1)(33) and tmr_registers(2)(33)) or                                                       
                            (tmr_registers(0)(33) and tmr_registers(2)(33));                                                         
                                                                                                                                     
        global_tmr_voter(2)(34)  <=    (tmr_registers(0)(34) and tmr_registers(1)(34)) or                                            
                            (tmr_registers(1)(34) and tmr_registers(2)(34)) or                                                       
                            (tmr_registers(0)(34) and tmr_registers(2)(34));                                                         
                                                                                                                                     
        global_tmr_voter(2)(35)  <=    (tmr_registers(0)(35) and tmr_registers(1)(35)) or                                            
                            (tmr_registers(1)(35) and tmr_registers(2)(35)) or                                                       
                            (tmr_registers(0)(35) and tmr_registers(2)(35));                                                         
                                                                                                                                     
        global_tmr_voter(2)(36)  <=    (tmr_registers(0)(36) and tmr_registers(1)(36)) or                                            
                            (tmr_registers(1)(36) and tmr_registers(2)(36)) or                                                       
                            (tmr_registers(0)(36) and tmr_registers(2)(36));                                                         
                                                                                                                                     
        global_tmr_voter(2)(37)  <=    (tmr_registers(0)(37) and tmr_registers(1)(37)) or                                            
                            (tmr_registers(1)(37) and tmr_registers(2)(37)) or                                                       
                            (tmr_registers(0)(37) and tmr_registers(2)(37));                                                         
                                                                                                                                     
        global_tmr_voter(2)(38)  <=    (tmr_registers(0)(38) and tmr_registers(1)(38)) or                                            
                            (tmr_registers(1)(38) and tmr_registers(2)(38)) or                                                       
                            (tmr_registers(0)(38) and tmr_registers(2)(38));                                                         
                                                                                                                                     
        global_tmr_voter(2)(39)  <=    (tmr_registers(0)(39) and tmr_registers(1)(39)) or                                            
                            (tmr_registers(1)(39) and tmr_registers(2)(39)) or                                                       
                            (tmr_registers(0)(39) and tmr_registers(2)(39));                                                         
                                                                                                                                     
        global_tmr_voter(2)(40)  <=    (tmr_registers(0)(40) and tmr_registers(1)(40)) or                                            
                            (tmr_registers(1)(40) and tmr_registers(2)(40)) or                                                       
                            (tmr_registers(0)(40) and tmr_registers(2)(40));                                                         
                                                                                                                                     
        global_tmr_voter(2)(41)  <=    (tmr_registers(0)(41) and tmr_registers(1)(41)) or                                            
                            (tmr_registers(1)(41) and tmr_registers(2)(41)) or                                                       
                            (tmr_registers(0)(41) and tmr_registers(2)(41));                                                         
                                                                                                                                     
        global_tmr_voter(2)(42)  <=    (tmr_registers(0)(42) and tmr_registers(1)(42)) or                                            
                            (tmr_registers(1)(42) and tmr_registers(2)(42)) or                                                       
                            (tmr_registers(0)(42) and tmr_registers(2)(42));                                                         
                                                                                                                                     
        global_tmr_voter(2)(43)  <=    (tmr_registers(0)(43) and tmr_registers(1)(43)) or                                            
                            (tmr_registers(1)(43) and tmr_registers(2)(43)) or                                                       
                            (tmr_registers(0)(43) and tmr_registers(2)(43));                                                         
                                                                                                                                     
        global_tmr_voter(2)(44)  <=    (tmr_registers(0)(44) and tmr_registers(1)(44)) or                                            
                            (tmr_registers(1)(44) and tmr_registers(2)(44)) or                                                       
                            (tmr_registers(0)(44) and tmr_registers(2)(44));                                                         
                                                                                                                                     
        global_tmr_voter(2)(45)  <=    (tmr_registers(0)(45) and tmr_registers(1)(45)) or                                            
                            (tmr_registers(1)(45) and tmr_registers(2)(45)) or                                                       
                            (tmr_registers(0)(45) and tmr_registers(2)(45));                                                         
                                                                                                                                     
        global_tmr_voter(2)(46)  <=    (tmr_registers(0)(46) and tmr_registers(1)(46)) or                                            
                            (tmr_registers(1)(46) and tmr_registers(2)(46)) or                                                       
                            (tmr_registers(0)(46) and tmr_registers(2)(46));                                                         
                                                                                                                                     
        global_tmr_voter(2)(47)  <=    (tmr_registers(0)(47) and tmr_registers(1)(47)) or                                            
                            (tmr_registers(1)(47) and tmr_registers(2)(47)) or                                                       
                            (tmr_registers(0)(47) and tmr_registers(2)(47));                                                         
                                                                                                                                     
        global_tmr_voter(2)(48)  <=    (tmr_registers(0)(48) and tmr_registers(1)(48)) or                                            
                            (tmr_registers(1)(48) and tmr_registers(2)(48)) or                                                       
                            (tmr_registers(0)(48) and tmr_registers(2)(48));                                                         
                                                                                                                                     
        global_tmr_voter(2)(49)  <=    (tmr_registers(0)(49) and tmr_registers(1)(49)) or                                            
                            (tmr_registers(1)(49) and tmr_registers(2)(49)) or                                                       
                            (tmr_registers(0)(49) and tmr_registers(2)(49));                                                         
                                                                                                                                     
        global_tmr_voter(2)(50)  <=    (tmr_registers(0)(50) and tmr_registers(1)(50)) or                                            
                            (tmr_registers(1)(50) and tmr_registers(2)(50)) or                                                       
                            (tmr_registers(0)(50) and tmr_registers(2)(50));                                                         
                                                                                                                                     
        global_tmr_voter(2)(51)  <=    (tmr_registers(0)(51) and tmr_registers(1)(51)) or                                            
                            (tmr_registers(1)(51) and tmr_registers(2)(51)) or                                                       
                            (tmr_registers(0)(51) and tmr_registers(2)(51));                                                         
                                                                                                                                     
        global_tmr_voter(2)(52)  <=    (tmr_registers(0)(52) and tmr_registers(1)(52)) or                                            
                            (tmr_registers(1)(52) and tmr_registers(2)(52)) or                                                       
                            (tmr_registers(0)(52) and tmr_registers(2)(52));                                                         
                                                                                                                                     
        global_tmr_voter(2)(53)  <=    (tmr_registers(0)(53) and tmr_registers(1)(53)) or                                            
                            (tmr_registers(1)(53) and tmr_registers(2)(53)) or                                                       
                            (tmr_registers(0)(53) and tmr_registers(2)(53));                                                         
                                                                                                                                     
        global_tmr_voter(2)(54)  <=    (tmr_registers(0)(54) and tmr_registers(1)(54)) or                                            
                            (tmr_registers(1)(54) and tmr_registers(2)(54)) or                                                       
                            (tmr_registers(0)(54) and tmr_registers(2)(54));                                                         
                                                                                                                                     
        global_tmr_voter(2)(55)  <=    (tmr_registers(0)(55) and tmr_registers(1)(55)) or                                            
                            (tmr_registers(1)(55) and tmr_registers(2)(55)) or                                                       
                            (tmr_registers(0)(55) and tmr_registers(2)(55));                                                         
                                                                                                                                     
        global_tmr_voter(2)(56)  <=    (tmr_registers(0)(56) and tmr_registers(1)(56)) or                                            
                            (tmr_registers(1)(56) and tmr_registers(2)(56)) or                                                       
                            (tmr_registers(0)(56) and tmr_registers(2)(56));                                                         
                                                                                                                                     
        global_tmr_voter(2)(57)  <=    (tmr_registers(0)(57) and tmr_registers(1)(57)) or                                            
                            (tmr_registers(1)(57) and tmr_registers(2)(57)) or                                                       
                            (tmr_registers(0)(57) and tmr_registers(2)(57));                                                         
                                                                                                                                     
        global_tmr_voter(2)(58)  <=    (tmr_registers(0)(58) and tmr_registers(1)(58)) or                                            
                            (tmr_registers(1)(58) and tmr_registers(2)(58)) or                                                       
                            (tmr_registers(0)(58) and tmr_registers(2)(58));                                                         
                                                                                                                                     
        global_tmr_voter(2)(59)  <=    (tmr_registers(0)(59) and tmr_registers(1)(59)) or                                            
                            (tmr_registers(1)(59) and tmr_registers(2)(59)) or                                                       
                            (tmr_registers(0)(59) and tmr_registers(2)(59));                                                         
                                                                                                                                     
        global_tmr_voter(2)(60)  <=    (tmr_registers(0)(60) and tmr_registers(1)(60)) or                                            
                            (tmr_registers(1)(60) and tmr_registers(2)(60)) or                                                       
                            (tmr_registers(0)(60) and tmr_registers(2)(60));                                                         
                                                                                                                                     
        global_tmr_voter(2)(61)  <=    (tmr_registers(0)(61) and tmr_registers(1)(61)) or                                            
                            (tmr_registers(1)(61) and tmr_registers(2)(61)) or                                                       
                            (tmr_registers(0)(61) and tmr_registers(2)(61));                                                         
                                                                                                                                     
        global_tmr_voter(2)(62)  <=    (tmr_registers(0)(62) and tmr_registers(1)(62)) or                                            
                            (tmr_registers(1)(62) and tmr_registers(2)(62)) or                                                       
                            (tmr_registers(0)(62) and tmr_registers(2)(62));                                                         
                                                                                                                                     
        global_tmr_voter(2)(63)  <=    (tmr_registers(0)(63) and tmr_registers(1)(63)) or                                            
                            (tmr_registers(1)(63) and tmr_registers(2)(63)) or                                                       
                            (tmr_registers(0)(63) and tmr_registers(2)(63));                                                         
                                                                                                                                     
        global_tmr_voter(2)(64)  <=    (tmr_registers(0)(64) and tmr_registers(1)(64)) or                                            
                            (tmr_registers(1)(64) and tmr_registers(2)(64)) or                                                       
                            (tmr_registers(0)(64) and tmr_registers(2)(64));                                                         
                                                                                                                                     
        global_tmr_voter(2)(65)  <=    (tmr_registers(0)(65) and tmr_registers(1)(65)) or                                            
                            (tmr_registers(1)(65) and tmr_registers(2)(65)) or                                                       
                            (tmr_registers(0)(65) and tmr_registers(2)(65));                                                         
                                                                                                                                     
        global_tmr_voter(2)(66)  <=    (tmr_registers(0)(66) and tmr_registers(1)(66)) or                                            
                            (tmr_registers(1)(66) and tmr_registers(2)(66)) or                                                       
                            (tmr_registers(0)(66) and tmr_registers(2)(66));                                                         
                                                                                                                                     
        global_tmr_voter(2)(67)  <=    (tmr_registers(0)(67) and tmr_registers(1)(67)) or                                            
                            (tmr_registers(1)(67) and tmr_registers(2)(67)) or                                                       
                            (tmr_registers(0)(67) and tmr_registers(2)(67));                                                         
                                                                                                                                     
        global_tmr_voter(2)(68)  <=    (tmr_registers(0)(68) and tmr_registers(1)(68)) or                                            
                            (tmr_registers(1)(68) and tmr_registers(2)(68)) or                                                       
                            (tmr_registers(0)(68) and tmr_registers(2)(68));                                                         
                                                                                                                                     
        global_tmr_voter(2)(69)  <=    (tmr_registers(0)(69) and tmr_registers(1)(69)) or                                            
                            (tmr_registers(1)(69) and tmr_registers(2)(69)) or                                                       
                            (tmr_registers(0)(69) and tmr_registers(2)(69));                                                         
                                                                                                                                     
        global_tmr_voter(2)(70)  <=    (tmr_registers(0)(70) and tmr_registers(1)(70)) or                                            
                            (tmr_registers(1)(70) and tmr_registers(2)(70)) or                                                       
                            (tmr_registers(0)(70) and tmr_registers(2)(70));                                                         
                                                                                                                                     
        global_tmr_voter(2)(71)  <=    (tmr_registers(0)(71) and tmr_registers(1)(71)) or                                            
                            (tmr_registers(1)(71) and tmr_registers(2)(71)) or                                                       
                            (tmr_registers(0)(71) and tmr_registers(2)(71));                                                         
                                                                                                                                     
        global_tmr_voter(2)(72)  <=    (tmr_registers(0)(72) and tmr_registers(1)(72)) or                                            
                            (tmr_registers(1)(72) and tmr_registers(2)(72)) or                                                       
                            (tmr_registers(0)(72) and tmr_registers(2)(72));                                                         
                                                                                                                                     
        global_tmr_voter(2)(73)  <=    (tmr_registers(0)(73) and tmr_registers(1)(73)) or                                            
                            (tmr_registers(1)(73) and tmr_registers(2)(73)) or                                                       
                            (tmr_registers(0)(73) and tmr_registers(2)(73));                                                         
                                                                                                                                     
        global_tmr_voter(2)(74)  <=    (tmr_registers(0)(74) and tmr_registers(1)(74)) or                                            
                            (tmr_registers(1)(74) and tmr_registers(2)(74)) or                                                       
                            (tmr_registers(0)(74) and tmr_registers(2)(74));                                                         
                                                                                                                                     
        global_tmr_voter(2)(75)  <=    (tmr_registers(0)(75) and tmr_registers(1)(75)) or                                            
                            (tmr_registers(1)(75) and tmr_registers(2)(75)) or                                                       
                            (tmr_registers(0)(75) and tmr_registers(2)(75));                                                         
                                                                                                                                     
        global_tmr_voter(2)(76)  <=    (tmr_registers(0)(76) and tmr_registers(1)(76)) or                                            
                            (tmr_registers(1)(76) and tmr_registers(2)(76)) or                                                       
                            (tmr_registers(0)(76) and tmr_registers(2)(76));                                                         
                                                                                                                                     
        global_tmr_voter(2)(77)  <=    (tmr_registers(0)(77) and tmr_registers(1)(77)) or                                            
                            (tmr_registers(1)(77) and tmr_registers(2)(77)) or                                                       
                            (tmr_registers(0)(77) and tmr_registers(2)(77));                                                         
                                                                                                                                     
        global_tmr_voter(2)(78)  <=    (tmr_registers(0)(78) and tmr_registers(1)(78)) or                                            
                            (tmr_registers(1)(78) and tmr_registers(2)(78)) or                                                       
                            (tmr_registers(0)(78) and tmr_registers(2)(78));                                                         
                                                                                                                                     
        global_tmr_voter(2)(79)  <=    (tmr_registers(0)(79) and tmr_registers(1)(79)) or                                            
                            (tmr_registers(1)(79) and tmr_registers(2)(79)) or                                                       
                            (tmr_registers(0)(79) and tmr_registers(2)(79));                                                         
                                                                                                                                     
        global_tmr_voter(2)(80)  <=    (tmr_registers(0)(80) and tmr_registers(1)(80)) or                                            
                            (tmr_registers(1)(80) and tmr_registers(2)(80)) or                                                       
                            (tmr_registers(0)(80) and tmr_registers(2)(80));                                                         
                                                                                                                                     
        global_tmr_voter(2)(81)  <=    (tmr_registers(0)(81) and tmr_registers(1)(81)) or                                            
                            (tmr_registers(1)(81) and tmr_registers(2)(81)) or                                                       
                            (tmr_registers(0)(81) and tmr_registers(2)(81));                                                         
                                                                                                                                     
        global_tmr_voter(2)(82)  <=    (tmr_registers(0)(82) and tmr_registers(1)(82)) or                                            
                            (tmr_registers(1)(82) and tmr_registers(2)(82)) or                                                       
                            (tmr_registers(0)(82) and tmr_registers(2)(82));                                                         
                                                                                                                                     
        global_tmr_voter(2)(83)  <=    (tmr_registers(0)(83) and tmr_registers(1)(83)) or                                            
                            (tmr_registers(1)(83) and tmr_registers(2)(83)) or                                                       
                            (tmr_registers(0)(83) and tmr_registers(2)(83));                                                         
                                                                                                                                     
        global_tmr_voter(2)(84)  <=    (tmr_registers(0)(84) and tmr_registers(1)(84)) or                                            
                            (tmr_registers(1)(84) and tmr_registers(2)(84)) or                                                       
                            (tmr_registers(0)(84) and tmr_registers(2)(84));                                                         
                                                                                                                                     
        global_tmr_voter(2)(85)  <=    (tmr_registers(0)(85) and tmr_registers(1)(85)) or                                            
                            (tmr_registers(1)(85) and tmr_registers(2)(85)) or                                                       
                            (tmr_registers(0)(85) and tmr_registers(2)(85));                                                         
                                                                                                                                     
        global_tmr_voter(2)(86)  <=    (tmr_registers(0)(86) and tmr_registers(1)(86)) or                                            
                            (tmr_registers(1)(86) and tmr_registers(2)(86)) or                                                       
                            (tmr_registers(0)(86) and tmr_registers(2)(86));                                                         
                                                                                                                                     
        global_tmr_voter(2)(87)  <=    (tmr_registers(0)(87) and tmr_registers(1)(87)) or                                            
                            (tmr_registers(1)(87) and tmr_registers(2)(87)) or                                                       
                            (tmr_registers(0)(87) and tmr_registers(2)(87));                                                         
                                                                                                                                     
        global_tmr_voter(2)(88)  <=    (tmr_registers(0)(88) and tmr_registers(1)(88)) or                                            
                            (tmr_registers(1)(88) and tmr_registers(2)(88)) or                                                       
                            (tmr_registers(0)(88) and tmr_registers(2)(88));                                                         
                                                                                                                                     
        global_tmr_voter(2)(89)  <=    (tmr_registers(0)(89) and tmr_registers(1)(89)) or                                            
                            (tmr_registers(1)(89) and tmr_registers(2)(89)) or                                                       
                            (tmr_registers(0)(89) and tmr_registers(2)(89));                                                         
                                                                                                                                     
        global_tmr_voter(2)(90)  <=    (tmr_registers(0)(90) and tmr_registers(1)(90)) or                                            
                            (tmr_registers(1)(90) and tmr_registers(2)(90)) or                                                       
                            (tmr_registers(0)(90) and tmr_registers(2)(90));                                                         
                                                                                                                                     
        global_tmr_voter(2)(91)  <=    (tmr_registers(0)(91) and tmr_registers(1)(91)) or                                            
                            (tmr_registers(1)(91) and tmr_registers(2)(91)) or                                                       
                            (tmr_registers(0)(91) and tmr_registers(2)(91));                                                         
                                                                                                                                     
        global_tmr_voter(2)(92)  <=    (tmr_registers(0)(92) and tmr_registers(1)(92)) or                                            
                            (tmr_registers(1)(92) and tmr_registers(2)(92)) or                                                       
                            (tmr_registers(0)(92) and tmr_registers(2)(92));                                                         
                                                                                                                                     
        global_tmr_voter(2)(93)  <=    (tmr_registers(0)(93) and tmr_registers(1)(93)) or                                            
                            (tmr_registers(1)(93) and tmr_registers(2)(93)) or                                                       
                            (tmr_registers(0)(93) and tmr_registers(2)(93));                                                         
                                                                                                                                     
        global_tmr_voter(2)(94)  <=    (tmr_registers(0)(94) and tmr_registers(1)(94)) or                                            
                            (tmr_registers(1)(94) and tmr_registers(2)(94)) or                                                       
                            (tmr_registers(0)(94) and tmr_registers(2)(94));                                                         
                                                                                                                                     
        global_tmr_voter(2)(95)  <=    (tmr_registers(0)(95) and tmr_registers(1)(95)) or                                            
                            (tmr_registers(1)(95) and tmr_registers(2)(95)) or                                                       
                            (tmr_registers(0)(95) and tmr_registers(2)(95));                                                         
                                                                                                                                     
        global_tmr_voter(2)(96)  <=    (tmr_registers(0)(96) and tmr_registers(1)(96)) or                                            
                            (tmr_registers(1)(96) and tmr_registers(2)(96)) or                                                       
                            (tmr_registers(0)(96) and tmr_registers(2)(96));                                                         
                                                                                                                                     
        global_tmr_voter(2)(97)  <=    (tmr_registers(0)(97) and tmr_registers(1)(97)) or                                            
                            (tmr_registers(1)(97) and tmr_registers(2)(97)) or                                                       
                            (tmr_registers(0)(97) and tmr_registers(2)(97));                                                         
                                                                                                                                     
        global_tmr_voter(2)(98)  <=    (tmr_registers(0)(98) and tmr_registers(1)(98)) or                                            
                            (tmr_registers(1)(98) and tmr_registers(2)(98)) or                                                       
                            (tmr_registers(0)(98) and tmr_registers(2)(98));                                                         
                                                                                                                                     
        global_tmr_voter(2)(99)  <=    (tmr_registers(0)(99) and tmr_registers(1)(99)) or                                            
                            (tmr_registers(1)(99) and tmr_registers(2)(99)) or                                                       
                            (tmr_registers(0)(99) and tmr_registers(2)(99));                                                         
                                                                                                                                     
        global_tmr_voter(2)(100)  <=    (tmr_registers(0)(100) and tmr_registers(1)(100)) or                                            
                            (tmr_registers(1)(100) and tmr_registers(2)(100)) or                                                       
                            (tmr_registers(0)(100) and tmr_registers(2)(100));                                                         
                                                                                                                                     
        global_tmr_voter(2)(101)  <=    (tmr_registers(0)(101) and tmr_registers(1)(101)) or                                            
                            (tmr_registers(1)(101) and tmr_registers(2)(101)) or                                                       
                            (tmr_registers(0)(101) and tmr_registers(2)(101));                                                         
                                                                                                                                     
        global_tmr_voter(2)(102)  <=    (tmr_registers(0)(102) and tmr_registers(1)(102)) or                                            
                            (tmr_registers(1)(102) and tmr_registers(2)(102)) or                                                       
                            (tmr_registers(0)(102) and tmr_registers(2)(102));                                                         
                                                                                                                                     
        global_tmr_voter(2)(103)  <=    (tmr_registers(0)(103) and tmr_registers(1)(103)) or                                            
                            (tmr_registers(1)(103) and tmr_registers(2)(103)) or                                                       
                            (tmr_registers(0)(103) and tmr_registers(2)(103));                                                         
                                                                                                                                     
        global_tmr_voter(2)(104)  <=    (tmr_registers(0)(104) and tmr_registers(1)(104)) or                                            
                            (tmr_registers(1)(104) and tmr_registers(2)(104)) or                                                       
                            (tmr_registers(0)(104) and tmr_registers(2)(104));                                                         
                                                                                                                                     
        global_tmr_voter(2)(105)  <=    (tmr_registers(0)(105) and tmr_registers(1)(105)) or                                            
                            (tmr_registers(1)(105) and tmr_registers(2)(105)) or                                                       
                            (tmr_registers(0)(105) and tmr_registers(2)(105));                                                         
                                                                                                                                     
        global_tmr_voter(2)(106)  <=    (tmr_registers(0)(106) and tmr_registers(1)(106)) or                                            
                            (tmr_registers(1)(106) and tmr_registers(2)(106)) or                                                       
                            (tmr_registers(0)(106) and tmr_registers(2)(106));                                                         
                                                                                                                                     
        global_tmr_voter(2)(107)  <=    (tmr_registers(0)(107) and tmr_registers(1)(107)) or                                            
                            (tmr_registers(1)(107) and tmr_registers(2)(107)) or                                                       
                            (tmr_registers(0)(107) and tmr_registers(2)(107));                                                         
                                                                                                                                     
        global_tmr_voter(2)(108)  <=    (tmr_registers(0)(108) and tmr_registers(1)(108)) or                                            
                            (tmr_registers(1)(108) and tmr_registers(2)(108)) or                                                       
                            (tmr_registers(0)(108) and tmr_registers(2)(108));                                                         
                                                                                                                                     
        global_tmr_voter(2)(109)  <=    (tmr_registers(0)(109) and tmr_registers(1)(109)) or                                            
                            (tmr_registers(1)(109) and tmr_registers(2)(109)) or                                                       
                            (tmr_registers(0)(109) and tmr_registers(2)(109));                                                         
                                                                                                                                     
        global_tmr_voter(2)(110)  <=    (tmr_registers(0)(110) and tmr_registers(1)(110)) or                                            
                            (tmr_registers(1)(110) and tmr_registers(2)(110)) or                                                       
                            (tmr_registers(0)(110) and tmr_registers(2)(110));                                                         
                                                                                                                                     
        global_tmr_voter(2)(111)  <=    (tmr_registers(0)(111) and tmr_registers(1)(111)) or                                            
                            (tmr_registers(1)(111) and tmr_registers(2)(111)) or                                                       
                            (tmr_registers(0)(111) and tmr_registers(2)(111));                                                         
                                                                                                                                     
        global_tmr_voter(2)(112)  <=    (tmr_registers(0)(112) and tmr_registers(1)(112)) or                                            
                            (tmr_registers(1)(112) and tmr_registers(2)(112)) or                                                       
                            (tmr_registers(0)(112) and tmr_registers(2)(112));                                                         
                                                                                                                                     
        global_tmr_voter(2)(113)  <=    (tmr_registers(0)(113) and tmr_registers(1)(113)) or                                            
                            (tmr_registers(1)(113) and tmr_registers(2)(113)) or                                                       
                            (tmr_registers(0)(113) and tmr_registers(2)(113));                                                         
                                                                                                                                     
        global_tmr_voter(2)(114)  <=    (tmr_registers(0)(114) and tmr_registers(1)(114)) or                                            
                            (tmr_registers(1)(114) and tmr_registers(2)(114)) or                                                       
                            (tmr_registers(0)(114) and tmr_registers(2)(114));                                                         
                                                                                                                                     
        global_tmr_voter(2)(115)  <=    (tmr_registers(0)(115) and tmr_registers(1)(115)) or                                            
                            (tmr_registers(1)(115) and tmr_registers(2)(115)) or                                                       
                            (tmr_registers(0)(115) and tmr_registers(2)(115));                                                         
                                                                                                                                     
        global_tmr_voter(2)(116)  <=    (tmr_registers(0)(116) and tmr_registers(1)(116)) or                                            
                            (tmr_registers(1)(116) and tmr_registers(2)(116)) or                                                       
                            (tmr_registers(0)(116) and tmr_registers(2)(116));                                                         
                                                                                                                                     
        global_tmr_voter(2)(117)  <=    (tmr_registers(0)(117) and tmr_registers(1)(117)) or                                            
                            (tmr_registers(1)(117) and tmr_registers(2)(117)) or                                                       
                            (tmr_registers(0)(117) and tmr_registers(2)(117));                                                         
                                                                                                                                     
        global_tmr_voter(2)(118)  <=    (tmr_registers(0)(118) and tmr_registers(1)(118)) or                                            
                            (tmr_registers(1)(118) and tmr_registers(2)(118)) or                                                       
                            (tmr_registers(0)(118) and tmr_registers(2)(118));                                                         
                                                                                                                                     
        global_tmr_voter(2)(119)  <=    (tmr_registers(0)(119) and tmr_registers(1)(119)) or                                            
                            (tmr_registers(1)(119) and tmr_registers(2)(119)) or                                                       
                            (tmr_registers(0)(119) and tmr_registers(2)(119));                                                         
                                                                                                                                     
        global_tmr_voter(2)(120)  <=    (tmr_registers(0)(120) and tmr_registers(1)(120)) or                                            
                            (tmr_registers(1)(120) and tmr_registers(2)(120)) or                                                       
                            (tmr_registers(0)(120) and tmr_registers(2)(120));                                                         
                                                                                                                                     
        global_tmr_voter(2)(121)  <=    (tmr_registers(0)(121) and tmr_registers(1)(121)) or                                            
                            (tmr_registers(1)(121) and tmr_registers(2)(121)) or                                                       
                            (tmr_registers(0)(121) and tmr_registers(2)(121));                                                         
                                                                                                                                     
        global_tmr_voter(2)(122)  <=    (tmr_registers(0)(122) and tmr_registers(1)(122)) or                                            
                            (tmr_registers(1)(122) and tmr_registers(2)(122)) or                                                       
                            (tmr_registers(0)(122) and tmr_registers(2)(122));                                                         
                                                                                                                                     
        global_tmr_voter(2)(123)  <=    (tmr_registers(0)(123) and tmr_registers(1)(123)) or                                            
                            (tmr_registers(1)(123) and tmr_registers(2)(123)) or                                                       
                            (tmr_registers(0)(123) and tmr_registers(2)(123));                                                         
                                                                                                                                     
        global_tmr_voter(2)(124)  <=    (tmr_registers(0)(124) and tmr_registers(1)(124)) or                                            
                            (tmr_registers(1)(124) and tmr_registers(2)(124)) or                                                       
                            (tmr_registers(0)(124) and tmr_registers(2)(124));                                                         
                                                                                                                                     
        global_tmr_voter(2)(125)  <=    (tmr_registers(0)(125) and tmr_registers(1)(125)) or                                            
                            (tmr_registers(1)(125) and tmr_registers(2)(125)) or                                                       
                            (tmr_registers(0)(125) and tmr_registers(2)(125));                                                         
                                                                                                                                     
        global_tmr_voter(2)(126)  <=    (tmr_registers(0)(126) and tmr_registers(1)(126)) or                                            
                            (tmr_registers(1)(126) and tmr_registers(2)(126)) or                                                       
                            (tmr_registers(0)(126) and tmr_registers(2)(126));                                                         
                                                                                                                                     
        global_tmr_voter(2)(127)  <=    (tmr_registers(0)(127) and tmr_registers(1)(127)) or                                            
                            (tmr_registers(1)(127) and tmr_registers(2)(127)) or                                                       
                            (tmr_registers(0)(127) and tmr_registers(2)(127));                                                         
                                                                                                                                     
        global_tmr_voter(2)(128)  <=    (tmr_registers(0)(128) and tmr_registers(1)(128)) or                                            
                            (tmr_registers(1)(128) and tmr_registers(2)(128)) or                                                       
                            (tmr_registers(0)(128) and tmr_registers(2)(128));                                                         
                                                                                                                                     
        global_tmr_voter(2)(129)  <=    (tmr_registers(0)(129) and tmr_registers(1)(129)) or                                            
                            (tmr_registers(1)(129) and tmr_registers(2)(129)) or                                                       
                            (tmr_registers(0)(129) and tmr_registers(2)(129));                                                         
                                                                                                                                     
        global_tmr_voter(2)(130)  <=    (tmr_registers(0)(130) and tmr_registers(1)(130)) or                                            
                            (tmr_registers(1)(130) and tmr_registers(2)(130)) or                                                       
                            (tmr_registers(0)(130) and tmr_registers(2)(130));                                                         
                                                                                                                                     
        global_tmr_voter(2)(131)  <=    (tmr_registers(0)(131) and tmr_registers(1)(131)) or                                            
                            (tmr_registers(1)(131) and tmr_registers(2)(131)) or                                                       
                            (tmr_registers(0)(131) and tmr_registers(2)(131));                                                         
                                                                                                                                     
        global_tmr_voter(2)(132)  <=    (tmr_registers(0)(132) and tmr_registers(1)(132)) or                                            
                            (tmr_registers(1)(132) and tmr_registers(2)(132)) or                                                       
                            (tmr_registers(0)(132) and tmr_registers(2)(132));                                                         
                                                                                                                                     
        global_tmr_voter(2)(133)  <=    (tmr_registers(0)(133) and tmr_registers(1)(133)) or                                            
                            (tmr_registers(1)(133) and tmr_registers(2)(133)) or                                                       
                            (tmr_registers(0)(133) and tmr_registers(2)(133));                                                         
                                                                                                                                     
        global_tmr_voter(2)(134)  <=    (tmr_registers(0)(134) and tmr_registers(1)(134)) or                                            
                            (tmr_registers(1)(134) and tmr_registers(2)(134)) or                                                       
                            (tmr_registers(0)(134) and tmr_registers(2)(134));                                                         
                                                                                                                                     
        global_tmr_voter(2)(135)  <=    (tmr_registers(0)(135) and tmr_registers(1)(135)) or                                            
                            (tmr_registers(1)(135) and tmr_registers(2)(135)) or                                                       
                            (tmr_registers(0)(135) and tmr_registers(2)(135));                                                         
                                                                                                                                     
        global_tmr_voter(2)(136)  <=    (tmr_registers(0)(136) and tmr_registers(1)(136)) or                                            
                            (tmr_registers(1)(136) and tmr_registers(2)(136)) or                                                       
                            (tmr_registers(0)(136) and tmr_registers(2)(136));                                                         
                                                                                                                                     
        global_tmr_voter(2)(137)  <=    (tmr_registers(0)(137) and tmr_registers(1)(137)) or                                            
                            (tmr_registers(1)(137) and tmr_registers(2)(137)) or                                                       
                            (tmr_registers(0)(137) and tmr_registers(2)(137));                                                         
                                                                                                                                     
        global_tmr_voter(2)(138)  <=    (tmr_registers(0)(138) and tmr_registers(1)(138)) or                                            
                            (tmr_registers(1)(138) and tmr_registers(2)(138)) or                                                       
                            (tmr_registers(0)(138) and tmr_registers(2)(138));                                                         
                                                                                                                                     
        global_tmr_voter(2)(139)  <=    (tmr_registers(0)(139) and tmr_registers(1)(139)) or                                            
                            (tmr_registers(1)(139) and tmr_registers(2)(139)) or                                                       
                            (tmr_registers(0)(139) and tmr_registers(2)(139));                                                         
                                                                                                                                     
        global_tmr_voter(2)(140)  <=    (tmr_registers(0)(140) and tmr_registers(1)(140)) or                                            
                            (tmr_registers(1)(140) and tmr_registers(2)(140)) or                                                       
                            (tmr_registers(0)(140) and tmr_registers(2)(140));                                                         
                                                                                                                                     
        global_tmr_voter(2)(141)  <=    (tmr_registers(0)(141) and tmr_registers(1)(141)) or                                            
                            (tmr_registers(1)(141) and tmr_registers(2)(141)) or                                                       
                            (tmr_registers(0)(141) and tmr_registers(2)(141));                                                         
                                                                                                                                     
        global_tmr_voter(2)(142)  <=    (tmr_registers(0)(142) and tmr_registers(1)(142)) or                                            
                            (tmr_registers(1)(142) and tmr_registers(2)(142)) or                                                       
                            (tmr_registers(0)(142) and tmr_registers(2)(142));                                                         
                                                                                                                                     
        global_tmr_voter(2)(143)  <=    (tmr_registers(0)(143) and tmr_registers(1)(143)) or                                            
                            (tmr_registers(1)(143) and tmr_registers(2)(143)) or                                                       
                            (tmr_registers(0)(143) and tmr_registers(2)(143));                                                         
                                                                                                                                     
        global_tmr_voter(2)(144)  <=    (tmr_registers(0)(144) and tmr_registers(1)(144)) or                                            
                            (tmr_registers(1)(144) and tmr_registers(2)(144)) or                                                       
                            (tmr_registers(0)(144) and tmr_registers(2)(144));                                                         
                                                                                                                                     
        global_tmr_voter(2)(145)  <=    (tmr_registers(0)(145) and tmr_registers(1)(145)) or                                            
                            (tmr_registers(1)(145) and tmr_registers(2)(145)) or                                                       
                            (tmr_registers(0)(145) and tmr_registers(2)(145));                                                         
                                                                                                                                     
        global_tmr_voter(2)(146)  <=    (tmr_registers(0)(146) and tmr_registers(1)(146)) or                                            
                            (tmr_registers(1)(146) and tmr_registers(2)(146)) or                                                       
                            (tmr_registers(0)(146) and tmr_registers(2)(146));                                                         
                                                                                                                                     
        global_tmr_voter(2)(147)  <=    (tmr_registers(0)(147) and tmr_registers(1)(147)) or                                            
                            (tmr_registers(1)(147) and tmr_registers(2)(147)) or                                                       
                            (tmr_registers(0)(147) and tmr_registers(2)(147));                                                         
                                                                                                                                     
        global_tmr_voter(2)(148)  <=    (tmr_registers(0)(148) and tmr_registers(1)(148)) or                                            
                            (tmr_registers(1)(148) and tmr_registers(2)(148)) or                                                       
                            (tmr_registers(0)(148) and tmr_registers(2)(148));                                                         
                                                                                                                                     
        global_tmr_voter(2)(149)  <=    (tmr_registers(0)(149) and tmr_registers(1)(149)) or                                            
                            (tmr_registers(1)(149) and tmr_registers(2)(149)) or                                                       
                            (tmr_registers(0)(149) and tmr_registers(2)(149));                                                         
                                                                                                                                     
        global_tmr_voter(2)(150)  <=    (tmr_registers(0)(150) and tmr_registers(1)(150)) or                                            
                            (tmr_registers(1)(150) and tmr_registers(2)(150)) or                                                       
                            (tmr_registers(0)(150) and tmr_registers(2)(150));                                                         
                                                                                                                                     
        global_tmr_voter(2)(151)  <=    (tmr_registers(0)(151) and tmr_registers(1)(151)) or                                            
                            (tmr_registers(1)(151) and tmr_registers(2)(151)) or                                                       
                            (tmr_registers(0)(151) and tmr_registers(2)(151));                                                         
                                                                                                                                     
        global_tmr_voter(2)(152)  <=    (tmr_registers(0)(152) and tmr_registers(1)(152)) or                                            
                            (tmr_registers(1)(152) and tmr_registers(2)(152)) or                                                       
                            (tmr_registers(0)(152) and tmr_registers(2)(152));                                                         
                                                                                                                                     
        global_tmr_voter(2)(153)  <=    (tmr_registers(0)(153) and tmr_registers(1)(153)) or                                            
                            (tmr_registers(1)(153) and tmr_registers(2)(153)) or                                                       
                            (tmr_registers(0)(153) and tmr_registers(2)(153));                                                         
                                                                                                                                     
        global_tmr_voter(2)(154)  <=    (tmr_registers(0)(154) and tmr_registers(1)(154)) or                                            
                            (tmr_registers(1)(154) and tmr_registers(2)(154)) or                                                       
                            (tmr_registers(0)(154) and tmr_registers(2)(154));                                                         
                                                                                                                                     
        global_tmr_voter(2)(155)  <=    (tmr_registers(0)(155) and tmr_registers(1)(155)) or                                            
                            (tmr_registers(1)(155) and tmr_registers(2)(155)) or                                                       
                            (tmr_registers(0)(155) and tmr_registers(2)(155));                                                         
                                                                                                                                     
        global_tmr_voter(2)(156)  <=    (tmr_registers(0)(156) and tmr_registers(1)(156)) or                                            
                            (tmr_registers(1)(156) and tmr_registers(2)(156)) or                                                       
                            (tmr_registers(0)(156) and tmr_registers(2)(156));                                                         
                                                                                                                                     
        global_tmr_voter(2)(157)  <=    (tmr_registers(0)(157) and tmr_registers(1)(157)) or                                            
                            (tmr_registers(1)(157) and tmr_registers(2)(157)) or                                                       
                            (tmr_registers(0)(157) and tmr_registers(2)(157));                                                         
                                                                                                                                     
        global_tmr_voter(2)(158)  <=    (tmr_registers(0)(158) and tmr_registers(1)(158)) or                                            
                            (tmr_registers(1)(158) and tmr_registers(2)(158)) or                                                       
                            (tmr_registers(0)(158) and tmr_registers(2)(158));                                                         
                                                                                                                                     
        global_tmr_voter(2)(159)  <=    (tmr_registers(0)(159) and tmr_registers(1)(159)) or                                            
                            (tmr_registers(1)(159) and tmr_registers(2)(159)) or                                                       
                            (tmr_registers(0)(159) and tmr_registers(2)(159));                                                         
                                                                                                                                     
        global_tmr_voter(2)(160)  <=    (tmr_registers(0)(160) and tmr_registers(1)(160)) or                                            
                            (tmr_registers(1)(160) and tmr_registers(2)(160)) or                                                       
                            (tmr_registers(0)(160) and tmr_registers(2)(160));                                                         
                                                                                                                                     
        global_tmr_voter(2)(161)  <=    (tmr_registers(0)(161) and tmr_registers(1)(161)) or                                            
                            (tmr_registers(1)(161) and tmr_registers(2)(161)) or                                                       
                            (tmr_registers(0)(161) and tmr_registers(2)(161));                                                         
                                                                                                                                     
        global_tmr_voter(2)(162)  <=    (tmr_registers(0)(162) and tmr_registers(1)(162)) or                                            
                            (tmr_registers(1)(162) and tmr_registers(2)(162)) or                                                       
                            (tmr_registers(0)(162) and tmr_registers(2)(162));                                                         
                                                                                                                                     
        global_tmr_voter(2)(163)  <=    (tmr_registers(0)(163) and tmr_registers(1)(163)) or                                            
                            (tmr_registers(1)(163) and tmr_registers(2)(163)) or                                                       
                            (tmr_registers(0)(163) and tmr_registers(2)(163));                                                         
                                                                                                                                     
        global_tmr_voter(2)(164)  <=    (tmr_registers(0)(164) and tmr_registers(1)(164)) or                                            
                            (tmr_registers(1)(164) and tmr_registers(2)(164)) or                                                       
                            (tmr_registers(0)(164) and tmr_registers(2)(164));                                                         
                                                                                                                                     
        global_tmr_voter(2)(165)  <=    (tmr_registers(0)(165) and tmr_registers(1)(165)) or                                            
                            (tmr_registers(1)(165) and tmr_registers(2)(165)) or                                                       
                            (tmr_registers(0)(165) and tmr_registers(2)(165));                                                         
                                                                                                                                     
        global_tmr_voter(2)(166)  <=    (tmr_registers(0)(166) and tmr_registers(1)(166)) or                                            
                            (tmr_registers(1)(166) and tmr_registers(2)(166)) or                                                       
                            (tmr_registers(0)(166) and tmr_registers(2)(166));                                                         
                                                                                                                                     
        global_tmr_voter(2)(167)  <=    (tmr_registers(0)(167) and tmr_registers(1)(167)) or                                            
                            (tmr_registers(1)(167) and tmr_registers(2)(167)) or                                                       
                            (tmr_registers(0)(167) and tmr_registers(2)(167));                                                         
                                                                                                                                     
        global_tmr_voter(2)(168)  <=    (tmr_registers(0)(168) and tmr_registers(1)(168)) or                                            
                            (tmr_registers(1)(168) and tmr_registers(2)(168)) or                                                       
                            (tmr_registers(0)(168) and tmr_registers(2)(168));                                                         
                                                                                                                                     
        global_tmr_voter(2)(169)  <=    (tmr_registers(0)(169) and tmr_registers(1)(169)) or                                            
                            (tmr_registers(1)(169) and tmr_registers(2)(169)) or                                                       
                            (tmr_registers(0)(169) and tmr_registers(2)(169));                                                         
                                                                                                                                     
        global_tmr_voter(2)(170)  <=    (tmr_registers(0)(170) and tmr_registers(1)(170)) or                                            
                            (tmr_registers(1)(170) and tmr_registers(2)(170)) or                                                       
                            (tmr_registers(0)(170) and tmr_registers(2)(170));                                                         
                                                                                                                                     
        global_tmr_voter(2)(171)  <=    (tmr_registers(0)(171) and tmr_registers(1)(171)) or                                            
                            (tmr_registers(1)(171) and tmr_registers(2)(171)) or                                                       
                            (tmr_registers(0)(171) and tmr_registers(2)(171));                                                         
                                                                                                                                     
        global_tmr_voter(2)(172)  <=    (tmr_registers(0)(172) and tmr_registers(1)(172)) or                                            
                            (tmr_registers(1)(172) and tmr_registers(2)(172)) or                                                       
                            (tmr_registers(0)(172) and tmr_registers(2)(172));                                                         
                                                                                                                                     
        global_tmr_voter(2)(173)  <=    (tmr_registers(0)(173) and tmr_registers(1)(173)) or                                            
                            (tmr_registers(1)(173) and tmr_registers(2)(173)) or                                                       
                            (tmr_registers(0)(173) and tmr_registers(2)(173));                                                         
                                                                                                                                     
        global_tmr_voter(2)(174)  <=    (tmr_registers(0)(174) and tmr_registers(1)(174)) or                                            
                            (tmr_registers(1)(174) and tmr_registers(2)(174)) or                                                       
                            (tmr_registers(0)(174) and tmr_registers(2)(174));                                                         
                                                                                                                                     
        global_tmr_voter(2)(175)  <=    (tmr_registers(0)(175) and tmr_registers(1)(175)) or                                            
                            (tmr_registers(1)(175) and tmr_registers(2)(175)) or                                                       
                            (tmr_registers(0)(175) and tmr_registers(2)(175));                                                         
                                                                                                                                     
        global_tmr_voter(2)(176)  <=    (tmr_registers(0)(176) and tmr_registers(1)(176)) or                                            
                            (tmr_registers(1)(176) and tmr_registers(2)(176)) or                                                       
                            (tmr_registers(0)(176) and tmr_registers(2)(176));                                                         
                                                                                                                                     
        global_tmr_voter(2)(177)  <=    (tmr_registers(0)(177) and tmr_registers(1)(177)) or                                            
                            (tmr_registers(1)(177) and tmr_registers(2)(177)) or                                                       
                            (tmr_registers(0)(177) and tmr_registers(2)(177));                                                         
                                                                                                                                     
        global_tmr_voter(2)(178)  <=    (tmr_registers(0)(178) and tmr_registers(1)(178)) or                                            
                            (tmr_registers(1)(178) and tmr_registers(2)(178)) or                                                       
                            (tmr_registers(0)(178) and tmr_registers(2)(178));                                                         
                                                                                                                                     
        global_tmr_voter(2)(179)  <=    (tmr_registers(0)(179) and tmr_registers(1)(179)) or                                            
                            (tmr_registers(1)(179) and tmr_registers(2)(179)) or                                                       
                            (tmr_registers(0)(179) and tmr_registers(2)(179));                                                         
                                                                                                                                     
        global_tmr_voter(2)(180)  <=    (tmr_registers(0)(180) and tmr_registers(1)(180)) or                                            
                            (tmr_registers(1)(180) and tmr_registers(2)(180)) or                                                       
                            (tmr_registers(0)(180) and tmr_registers(2)(180));                                                         
                                                                                                                                     
        global_tmr_voter(2)(181)  <=    (tmr_registers(0)(181) and tmr_registers(1)(181)) or                                            
                            (tmr_registers(1)(181) and tmr_registers(2)(181)) or                                                       
                            (tmr_registers(0)(181) and tmr_registers(2)(181));                                                         
                                                                                                                                     
        global_tmr_voter(2)(182)  <=    (tmr_registers(0)(182) and tmr_registers(1)(182)) or                                            
                            (tmr_registers(1)(182) and tmr_registers(2)(182)) or                                                       
                            (tmr_registers(0)(182) and tmr_registers(2)(182));                                                         
                                                                                                                                     
        global_tmr_voter(2)(183)  <=    (tmr_registers(0)(183) and tmr_registers(1)(183)) or                                            
                            (tmr_registers(1)(183) and tmr_registers(2)(183)) or                                                       
                            (tmr_registers(0)(183) and tmr_registers(2)(183));                                                         
                                                                                                                                     
        global_tmr_voter(2)(184)  <=    (tmr_registers(0)(184) and tmr_registers(1)(184)) or                                            
                            (tmr_registers(1)(184) and tmr_registers(2)(184)) or                                                       
                            (tmr_registers(0)(184) and tmr_registers(2)(184));                                                         
                                                                                                                                     
        global_tmr_voter(2)(185)  <=    (tmr_registers(0)(185) and tmr_registers(1)(185)) or                                            
                            (tmr_registers(1)(185) and tmr_registers(2)(185)) or                                                       
                            (tmr_registers(0)(185) and tmr_registers(2)(185));                                                         
                                                                                                                                     
        global_tmr_voter(2)(186)  <=    (tmr_registers(0)(186) and tmr_registers(1)(186)) or                                            
                            (tmr_registers(1)(186) and tmr_registers(2)(186)) or                                                       
                            (tmr_registers(0)(186) and tmr_registers(2)(186));                                                         
                                                                                                                                     
        global_tmr_voter(2)(187)  <=    (tmr_registers(0)(187) and tmr_registers(1)(187)) or                                            
                            (tmr_registers(1)(187) and tmr_registers(2)(187)) or                                                       
                            (tmr_registers(0)(187) and tmr_registers(2)(187));                                                         
                                                                                                                                     
        global_tmr_voter(2)(188)  <=    (tmr_registers(0)(188) and tmr_registers(1)(188)) or                                            
                            (tmr_registers(1)(188) and tmr_registers(2)(188)) or                                                       
                            (tmr_registers(0)(188) and tmr_registers(2)(188));                                                         
                                                                                                                                     
        global_tmr_voter(2)(189)  <=    (tmr_registers(0)(189) and tmr_registers(1)(189)) or                                            
                            (tmr_registers(1)(189) and tmr_registers(2)(189)) or                                                       
                            (tmr_registers(0)(189) and tmr_registers(2)(189));                                                         
                                                                                                                                     
        global_tmr_voter(2)(190)  <=    (tmr_registers(0)(190) and tmr_registers(1)(190)) or                                            
                            (tmr_registers(1)(190) and tmr_registers(2)(190)) or                                                       
                            (tmr_registers(0)(190) and tmr_registers(2)(190));                                                         
                                                                                                                                     
        global_tmr_voter(2)(191)  <=    (tmr_registers(0)(191) and tmr_registers(1)(191)) or                                            
                            (tmr_registers(1)(191) and tmr_registers(2)(191)) or                                                       
                            (tmr_registers(0)(191) and tmr_registers(2)(191));                                                         
                                                                                                                                     
        global_tmr_voter(2)(192)  <=    (tmr_registers(0)(192) and tmr_registers(1)(192)) or                                            
                            (tmr_registers(1)(192) and tmr_registers(2)(192)) or                                                       
                            (tmr_registers(0)(192) and tmr_registers(2)(192));                                                         
                                                                                                                                     
        global_tmr_voter(2)(193)  <=    (tmr_registers(0)(193) and tmr_registers(1)(193)) or                                            
                            (tmr_registers(1)(193) and tmr_registers(2)(193)) or                                                       
                            (tmr_registers(0)(193) and tmr_registers(2)(193));                                                         
                                                                                                                                     
        global_tmr_voter(2)(194)  <=    (tmr_registers(0)(194) and tmr_registers(1)(194)) or                                            
                            (tmr_registers(1)(194) and tmr_registers(2)(194)) or                                                       
                            (tmr_registers(0)(194) and tmr_registers(2)(194));                                                         
                                                                                                                                     
        global_tmr_voter(2)(195)  <=    (tmr_registers(0)(195) and tmr_registers(1)(195)) or                                            
                            (tmr_registers(1)(195) and tmr_registers(2)(195)) or                                                       
                            (tmr_registers(0)(195) and tmr_registers(2)(195));                                                         
                                                                                                                                     
        global_tmr_voter(2)(196)  <=    (tmr_registers(0)(196) and tmr_registers(1)(196)) or                                            
                            (tmr_registers(1)(196) and tmr_registers(2)(196)) or                                                       
                            (tmr_registers(0)(196) and tmr_registers(2)(196));                                                         
                                                                                                                                     
        global_tmr_voter(2)(197)  <=    (tmr_registers(0)(197) and tmr_registers(1)(197)) or                                            
                            (tmr_registers(1)(197) and tmr_registers(2)(197)) or                                                       
                            (tmr_registers(0)(197) and tmr_registers(2)(197));                                                         
                                                                                                                                     
        global_tmr_voter(2)(198)  <=    (tmr_registers(0)(198) and tmr_registers(1)(198)) or                                            
                            (tmr_registers(1)(198) and tmr_registers(2)(198)) or                                                       
                            (tmr_registers(0)(198) and tmr_registers(2)(198));                                                         
                                                                                                                                     
        global_tmr_voter(2)(199)  <=    (tmr_registers(0)(199) and tmr_registers(1)(199)) or                                            
                            (tmr_registers(1)(199) and tmr_registers(2)(199)) or                                                       
                            (tmr_registers(0)(199) and tmr_registers(2)(199));                                                         
                                                                                                                                     
        global_tmr_voter(2)(200)  <=    (tmr_registers(0)(200) and tmr_registers(1)(200)) or                                            
                            (tmr_registers(1)(200) and tmr_registers(2)(200)) or                                                       
                            (tmr_registers(0)(200) and tmr_registers(2)(200));                                                         
                                                                                                                                     
        global_tmr_voter(2)(201)  <=    (tmr_registers(0)(201) and tmr_registers(1)(201)) or                                            
                            (tmr_registers(1)(201) and tmr_registers(2)(201)) or                                                       
                            (tmr_registers(0)(201) and tmr_registers(2)(201));                                                         
                                                                                                                                     
        global_tmr_voter(2)(202)  <=    (tmr_registers(0)(202) and tmr_registers(1)(202)) or                                            
                            (tmr_registers(1)(202) and tmr_registers(2)(202)) or                                                       
                            (tmr_registers(0)(202) and tmr_registers(2)(202));                                                         
                                                                                                                                     
        global_tmr_voter(2)(203)  <=    (tmr_registers(0)(203) and tmr_registers(1)(203)) or                                            
                            (tmr_registers(1)(203) and tmr_registers(2)(203)) or                                                       
                            (tmr_registers(0)(203) and tmr_registers(2)(203));                                                         
                                                                                                                                     
        global_tmr_voter(2)(204)  <=    (tmr_registers(0)(204) and tmr_registers(1)(204)) or                                            
                            (tmr_registers(1)(204) and tmr_registers(2)(204)) or                                                       
                            (tmr_registers(0)(204) and tmr_registers(2)(204));                                                         
                                                                                                                                     
        global_tmr_voter(2)(205)  <=    (tmr_registers(0)(205) and tmr_registers(1)(205)) or                                            
                            (tmr_registers(1)(205) and tmr_registers(2)(205)) or                                                       
                            (tmr_registers(0)(205) and tmr_registers(2)(205));                                                         
                                                                                                                                     
        global_tmr_voter(2)(206)  <=    (tmr_registers(0)(206) and tmr_registers(1)(206)) or                                            
                            (tmr_registers(1)(206) and tmr_registers(2)(206)) or                                                       
                            (tmr_registers(0)(206) and tmr_registers(2)(206));                                                         
                                                                                                                                     
        global_tmr_voter(2)(207)  <=    (tmr_registers(0)(207) and tmr_registers(1)(207)) or                                            
                            (tmr_registers(1)(207) and tmr_registers(2)(207)) or                                                       
                            (tmr_registers(0)(207) and tmr_registers(2)(207));                                                         
                                                                                                                                     
        global_tmr_voter(2)(208)  <=    (tmr_registers(0)(208) and tmr_registers(1)(208)) or                                            
                            (tmr_registers(1)(208) and tmr_registers(2)(208)) or                                                       
                            (tmr_registers(0)(208) and tmr_registers(2)(208));                                                         
                                                                                                                                     
        global_tmr_voter(2)(209)  <=    (tmr_registers(0)(209) and tmr_registers(1)(209)) or                                            
                            (tmr_registers(1)(209) and tmr_registers(2)(209)) or                                                       
                            (tmr_registers(0)(209) and tmr_registers(2)(209));                                                         
                                                                                                                                     
        global_tmr_voter(2)(210)  <=    (tmr_registers(0)(210) and tmr_registers(1)(210)) or                                            
                            (tmr_registers(1)(210) and tmr_registers(2)(210)) or                                                       
                            (tmr_registers(0)(210) and tmr_registers(2)(210));                                                         
                                                                                                                                     
        global_tmr_voter(2)(211)  <=    (tmr_registers(0)(211) and tmr_registers(1)(211)) or                                            
                            (tmr_registers(1)(211) and tmr_registers(2)(211)) or                                                       
                            (tmr_registers(0)(211) and tmr_registers(2)(211));                                                         
                                                                                                                                     
        global_tmr_voter(2)(212)  <=    (tmr_registers(0)(212) and tmr_registers(1)(212)) or                                            
                            (tmr_registers(1)(212) and tmr_registers(2)(212)) or                                                       
                            (tmr_registers(0)(212) and tmr_registers(2)(212));                                                         
                                                                                                                                     
        global_tmr_voter(2)(213)  <=    (tmr_registers(0)(213) and tmr_registers(1)(213)) or                                            
                            (tmr_registers(1)(213) and tmr_registers(2)(213)) or                                                       
                            (tmr_registers(0)(213) and tmr_registers(2)(213));                                                         
                                                                                                                                     
        global_tmr_voter(2)(214)  <=    (tmr_registers(0)(214) and tmr_registers(1)(214)) or                                            
                            (tmr_registers(1)(214) and tmr_registers(2)(214)) or                                                       
                            (tmr_registers(0)(214) and tmr_registers(2)(214));                                                         
                                                                                                                                     
        global_tmr_voter(2)(215)  <=    (tmr_registers(0)(215) and tmr_registers(1)(215)) or                                            
                            (tmr_registers(1)(215) and tmr_registers(2)(215)) or                                                       
                            (tmr_registers(0)(215) and tmr_registers(2)(215));                                                         
                                                                                                                                     
        global_tmr_voter(2)(216)  <=    (tmr_registers(0)(216) and tmr_registers(1)(216)) or                                            
                            (tmr_registers(1)(216) and tmr_registers(2)(216)) or                                                       
                            (tmr_registers(0)(216) and tmr_registers(2)(216));                                                         
                                                                                                                                     
        global_tmr_voter(2)(217)  <=    (tmr_registers(0)(217) and tmr_registers(1)(217)) or                                            
                            (tmr_registers(1)(217) and tmr_registers(2)(217)) or                                                       
                            (tmr_registers(0)(217) and tmr_registers(2)(217));                                                         
                                                                                                                                     
        global_tmr_voter(2)(218)  <=    (tmr_registers(0)(218) and tmr_registers(1)(218)) or                                            
                            (tmr_registers(1)(218) and tmr_registers(2)(218)) or                                                       
                            (tmr_registers(0)(218) and tmr_registers(2)(218));                                                         
                                                                                                                                     
        global_tmr_voter(2)(219)  <=    (tmr_registers(0)(219) and tmr_registers(1)(219)) or                                            
                            (tmr_registers(1)(219) and tmr_registers(2)(219)) or                                                       
                            (tmr_registers(0)(219) and tmr_registers(2)(219));                                                         
                                                                                                                                     
        global_tmr_voter(2)(220)  <=    (tmr_registers(0)(220) and tmr_registers(1)(220)) or                                            
                            (tmr_registers(1)(220) and tmr_registers(2)(220)) or                                                       
                            (tmr_registers(0)(220) and tmr_registers(2)(220));                                                         
                                                                                                                                     
        global_tmr_voter(2)(221)  <=    (tmr_registers(0)(221) and tmr_registers(1)(221)) or                                            
                            (tmr_registers(1)(221) and tmr_registers(2)(221)) or                                                       
                            (tmr_registers(0)(221) and tmr_registers(2)(221));                                                         
                                                                                                                                     
        global_tmr_voter(2)(222)  <=    (tmr_registers(0)(222) and tmr_registers(1)(222)) or                                            
                            (tmr_registers(1)(222) and tmr_registers(2)(222)) or                                                       
                            (tmr_registers(0)(222) and tmr_registers(2)(222));                                                         
                                                                                                                                     
        global_tmr_voter(2)(223)  <=    (tmr_registers(0)(223) and tmr_registers(1)(223)) or                                            
                            (tmr_registers(1)(223) and tmr_registers(2)(223)) or                                                       
                            (tmr_registers(0)(223) and tmr_registers(2)(223));                                                         
                                                                                                                                     
        global_tmr_voter(2)(224)  <=    (tmr_registers(0)(224) and tmr_registers(1)(224)) or                                            
                            (tmr_registers(1)(224) and tmr_registers(2)(224)) or                                                       
                            (tmr_registers(0)(224) and tmr_registers(2)(224));                                                         
                                                                                                                                     
        global_tmr_voter(2)(225)  <=    (tmr_registers(0)(225) and tmr_registers(1)(225)) or                                            
                            (tmr_registers(1)(225) and tmr_registers(2)(225)) or                                                       
                            (tmr_registers(0)(225) and tmr_registers(2)(225));                                                         
                                                                                                                                     
        global_tmr_voter(2)(226)  <=    (tmr_registers(0)(226) and tmr_registers(1)(226)) or                                            
                            (tmr_registers(1)(226) and tmr_registers(2)(226)) or                                                       
                            (tmr_registers(0)(226) and tmr_registers(2)(226));                                                         
                                                                                                                                     
        global_tmr_voter(2)(227)  <=    (tmr_registers(0)(227) and tmr_registers(1)(227)) or                                            
                            (tmr_registers(1)(227) and tmr_registers(2)(227)) or                                                       
                            (tmr_registers(0)(227) and tmr_registers(2)(227));                                                         
                                                                                                                                     
        global_tmr_voter(2)(228)  <=    (tmr_registers(0)(228) and tmr_registers(1)(228)) or                                            
                            (tmr_registers(1)(228) and tmr_registers(2)(228)) or                                                       
                            (tmr_registers(0)(228) and tmr_registers(2)(228));                                                         
                                                                                                                                     
        global_tmr_voter(2)(229)  <=    (tmr_registers(0)(229) and tmr_registers(1)(229)) or                                            
                            (tmr_registers(1)(229) and tmr_registers(2)(229)) or                                                       
                            (tmr_registers(0)(229) and tmr_registers(2)(229));                                                         
                                                                                                                                     
        global_tmr_voter(2)(230)  <=    (tmr_registers(0)(230) and tmr_registers(1)(230)) or                                            
                            (tmr_registers(1)(230) and tmr_registers(2)(230)) or                                                       
                            (tmr_registers(0)(230) and tmr_registers(2)(230));                                                         
                                                                                                                                     
        global_tmr_voter(2)(231)  <=    (tmr_registers(0)(231) and tmr_registers(1)(231)) or                                            
                            (tmr_registers(1)(231) and tmr_registers(2)(231)) or                                                       
                            (tmr_registers(0)(231) and tmr_registers(2)(231));                                                         
                                                                                                                                     
        global_tmr_voter(2)(232)  <=    (tmr_registers(0)(232) and tmr_registers(1)(232)) or                                            
                            (tmr_registers(1)(232) and tmr_registers(2)(232)) or                                                       
                            (tmr_registers(0)(232) and tmr_registers(2)(232));                                                         
                                                                                                                                     
        global_tmr_voter(2)(233)  <=    (tmr_registers(0)(233) and tmr_registers(1)(233)) or                                            
                            (tmr_registers(1)(233) and tmr_registers(2)(233)) or                                                       
                            (tmr_registers(0)(233) and tmr_registers(2)(233));                                                         
                                                                                                                                     
        global_tmr_voter(2)(234)  <=    (tmr_registers(0)(234) and tmr_registers(1)(234)) or                                            
                            (tmr_registers(1)(234) and tmr_registers(2)(234)) or                                                       
                            (tmr_registers(0)(234) and tmr_registers(2)(234));                                                         
                                                                                                                                     
        global_tmr_voter(2)(235)  <=    (tmr_registers(0)(235) and tmr_registers(1)(235)) or                                            
                            (tmr_registers(1)(235) and tmr_registers(2)(235)) or                                                       
                            (tmr_registers(0)(235) and tmr_registers(2)(235));                                                         
                                                                                                                                     
        global_tmr_voter(2)(236)  <=    (tmr_registers(0)(236) and tmr_registers(1)(236)) or                                            
                            (tmr_registers(1)(236) and tmr_registers(2)(236)) or                                                       
                            (tmr_registers(0)(236) and tmr_registers(2)(236));                                                         
                                                                                                                                     
        global_tmr_voter(2)(237)  <=    (tmr_registers(0)(237) and tmr_registers(1)(237)) or                                            
                            (tmr_registers(1)(237) and tmr_registers(2)(237)) or                                                       
                            (tmr_registers(0)(237) and tmr_registers(2)(237));                                                         
                                                                                                                                     
        global_tmr_voter(2)(238)  <=    (tmr_registers(0)(238) and tmr_registers(1)(238)) or                                            
                            (tmr_registers(1)(238) and tmr_registers(2)(238)) or                                                       
                            (tmr_registers(0)(238) and tmr_registers(2)(238));                                                         
                                                                                                                                     
        global_tmr_voter(2)(239)  <=    (tmr_registers(0)(239) and tmr_registers(1)(239)) or                                            
                            (tmr_registers(1)(239) and tmr_registers(2)(239)) or                                                       
                            (tmr_registers(0)(239) and tmr_registers(2)(239));                                                         
                                                                                                                                     
        global_tmr_voter(2)(240)  <=    (tmr_registers(0)(240) and tmr_registers(1)(240)) or                                            
                            (tmr_registers(1)(240) and tmr_registers(2)(240)) or                                                       
                            (tmr_registers(0)(240) and tmr_registers(2)(240));                                                         
                                                                                                                                     
        global_tmr_voter(2)(241)  <=    (tmr_registers(0)(241) and tmr_registers(1)(241)) or                                            
                            (tmr_registers(1)(241) and tmr_registers(2)(241)) or                                                       
                            (tmr_registers(0)(241) and tmr_registers(2)(241));                                                         
                                                                                                                                     
        global_tmr_voter(2)(242)  <=    (tmr_registers(0)(242) and tmr_registers(1)(242)) or                                            
                            (tmr_registers(1)(242) and tmr_registers(2)(242)) or                                                       
                            (tmr_registers(0)(242) and tmr_registers(2)(242));                                                         
                                                                                                                                     
        global_tmr_voter(2)(243)  <=    (tmr_registers(0)(243) and tmr_registers(1)(243)) or                                            
                            (tmr_registers(1)(243) and tmr_registers(2)(243)) or                                                       
                            (tmr_registers(0)(243) and tmr_registers(2)(243));                                                         
                                                                                                                                     
        global_tmr_voter(2)(244)  <=    (tmr_registers(0)(244) and tmr_registers(1)(244)) or                                            
                            (tmr_registers(1)(244) and tmr_registers(2)(244)) or                                                       
                            (tmr_registers(0)(244) and tmr_registers(2)(244));                                                         
                                                                                                                                     
        global_tmr_voter(2)(245)  <=    (tmr_registers(0)(245) and tmr_registers(1)(245)) or                                            
                            (tmr_registers(1)(245) and tmr_registers(2)(245)) or                                                       
                            (tmr_registers(0)(245) and tmr_registers(2)(245));                                                         
                                                                                                                                     
        global_tmr_voter(2)(246)  <=    (tmr_registers(0)(246) and tmr_registers(1)(246)) or                                            
                            (tmr_registers(1)(246) and tmr_registers(2)(246)) or                                                       
                            (tmr_registers(0)(246) and tmr_registers(2)(246));                                                         
                                                                                                                                     
        global_tmr_voter(2)(247)  <=    (tmr_registers(0)(247) and tmr_registers(1)(247)) or                                            
                            (tmr_registers(1)(247) and tmr_registers(2)(247)) or                                                       
                            (tmr_registers(0)(247) and tmr_registers(2)(247));                                                         
                                                                                                                                     
        global_tmr_voter(2)(248)  <=    (tmr_registers(0)(248) and tmr_registers(1)(248)) or                                            
                            (tmr_registers(1)(248) and tmr_registers(2)(248)) or                                                       
                            (tmr_registers(0)(248) and tmr_registers(2)(248));                                                         
                                                                                                                                     
        global_tmr_voter(2)(249)  <=    (tmr_registers(0)(249) and tmr_registers(1)(249)) or                                            
                            (tmr_registers(1)(249) and tmr_registers(2)(249)) or                                                       
                            (tmr_registers(0)(249) and tmr_registers(2)(249));                                                         
                                                                                                                                     
        global_tmr_voter(2)(250)  <=    (tmr_registers(0)(250) and tmr_registers(1)(250)) or                                            
                            (tmr_registers(1)(250) and tmr_registers(2)(250)) or                                                       
                            (tmr_registers(0)(250) and tmr_registers(2)(250));                                                         
                                                                                                                                     
        global_tmr_voter(2)(251)  <=    (tmr_registers(0)(251) and tmr_registers(1)(251)) or                                            
                            (tmr_registers(1)(251) and tmr_registers(2)(251)) or                                                       
                            (tmr_registers(0)(251) and tmr_registers(2)(251));                                                         
                                                                                                                                     
        global_tmr_voter(2)(252)  <=    (tmr_registers(0)(252) and tmr_registers(1)(252)) or                                            
                            (tmr_registers(1)(252) and tmr_registers(2)(252)) or                                                       
                            (tmr_registers(0)(252) and tmr_registers(2)(252));                                                         
                                                                                                                                     
        global_tmr_voter(2)(253)  <=    (tmr_registers(0)(253) and tmr_registers(1)(253)) or                                            
                            (tmr_registers(1)(253) and tmr_registers(2)(253)) or                                                       
                            (tmr_registers(0)(253) and tmr_registers(2)(253));                                                         
                                                                                                                                     
        global_tmr_voter(2)(254)  <=    (tmr_registers(0)(254) and tmr_registers(1)(254)) or                                            
                            (tmr_registers(1)(254) and tmr_registers(2)(254)) or                                                       
                            (tmr_registers(0)(254) and tmr_registers(2)(254));                                                         
                                                                                                                                     
        global_tmr_voter(2)(255)  <=    (tmr_registers(0)(255) and tmr_registers(1)(255)) or                                            
                            (tmr_registers(1)(255) and tmr_registers(2)(255)) or                                                       
                            (tmr_registers(0)(255) and tmr_registers(2)(255));                                                         
                                                                                                                                     
        global_tmr_voter(2)(256)  <=    (tmr_registers(0)(256) and tmr_registers(1)(256)) or                                            
                            (tmr_registers(1)(256) and tmr_registers(2)(256)) or                                                       
                            (tmr_registers(0)(256) and tmr_registers(2)(256));                                                         
                                                                                                                                     
        global_tmr_voter(2)(257)  <=    (tmr_registers(0)(257) and tmr_registers(1)(257)) or                                            
                            (tmr_registers(1)(257) and tmr_registers(2)(257)) or                                                       
                            (tmr_registers(0)(257) and tmr_registers(2)(257));                                                         
                                                                                                                                     
        global_tmr_voter(2)(258)  <=    (tmr_registers(0)(258) and tmr_registers(1)(258)) or                                            
                            (tmr_registers(1)(258) and tmr_registers(2)(258)) or                                                       
                            (tmr_registers(0)(258) and tmr_registers(2)(258));                                                         
                                                                                                                                     
        global_tmr_voter(2)(259)  <=    (tmr_registers(0)(259) and tmr_registers(1)(259)) or                                            
                            (tmr_registers(1)(259) and tmr_registers(2)(259)) or                                                       
                            (tmr_registers(0)(259) and tmr_registers(2)(259));                                                         
                                                                                                                                     
        global_tmr_voter(2)(260)  <=    (tmr_registers(0)(260) and tmr_registers(1)(260)) or                                            
                            (tmr_registers(1)(260) and tmr_registers(2)(260)) or                                                       
                            (tmr_registers(0)(260) and tmr_registers(2)(260));                                                         
                                                                                                                                     
        global_tmr_voter(2)(261)  <=    (tmr_registers(0)(261) and tmr_registers(1)(261)) or                                            
                            (tmr_registers(1)(261) and tmr_registers(2)(261)) or                                                       
                            (tmr_registers(0)(261) and tmr_registers(2)(261));                                                         
                                                                                                                                     
        global_tmr_voter(2)(262)  <=    (tmr_registers(0)(262) and tmr_registers(1)(262)) or                                            
                            (tmr_registers(1)(262) and tmr_registers(2)(262)) or                                                       
                            (tmr_registers(0)(262) and tmr_registers(2)(262));                                                         
                                                                                                                                     
        global_tmr_voter(2)(263)  <=    (tmr_registers(0)(263) and tmr_registers(1)(263)) or                                            
                            (tmr_registers(1)(263) and tmr_registers(2)(263)) or                                                       
                            (tmr_registers(0)(263) and tmr_registers(2)(263));                                                         
                                                                                                                                     
        global_tmr_voter(2)(264)  <=    (tmr_registers(0)(264) and tmr_registers(1)(264)) or                                            
                            (tmr_registers(1)(264) and tmr_registers(2)(264)) or                                                       
                            (tmr_registers(0)(264) and tmr_registers(2)(264));                                                         
                                                                                                                                     
        global_tmr_voter(2)(265)  <=    (tmr_registers(0)(265) and tmr_registers(1)(265)) or                                            
                            (tmr_registers(1)(265) and tmr_registers(2)(265)) or                                                       
                            (tmr_registers(0)(265) and tmr_registers(2)(265));                                                         
                                                                                                                                     
        global_tmr_voter(2)(266)  <=    (tmr_registers(0)(266) and tmr_registers(1)(266)) or                                            
                            (tmr_registers(1)(266) and tmr_registers(2)(266)) or                                                       
                            (tmr_registers(0)(266) and tmr_registers(2)(266));                                                         
                                                                                                                                     
        global_tmr_voter(2)(267)  <=    (tmr_registers(0)(267) and tmr_registers(1)(267)) or                                            
                            (tmr_registers(1)(267) and tmr_registers(2)(267)) or                                                       
                            (tmr_registers(0)(267) and tmr_registers(2)(267));                                                         
                                                                                                                                     
        global_tmr_voter(2)(268)  <=    (tmr_registers(0)(268) and tmr_registers(1)(268)) or                                            
                            (tmr_registers(1)(268) and tmr_registers(2)(268)) or                                                       
                            (tmr_registers(0)(268) and tmr_registers(2)(268));                                                         
                                                                                                                                     
        global_tmr_voter(2)(269)  <=    (tmr_registers(0)(269) and tmr_registers(1)(269)) or                                            
                            (tmr_registers(1)(269) and tmr_registers(2)(269)) or                                                       
                            (tmr_registers(0)(269) and tmr_registers(2)(269));                                                         
                                                                                                                                     
        global_tmr_voter(2)(270)  <=    (tmr_registers(0)(270) and tmr_registers(1)(270)) or                                            
                            (tmr_registers(1)(270) and tmr_registers(2)(270)) or                                                       
                            (tmr_registers(0)(270) and tmr_registers(2)(270));                                                         
                                                                                                                                     
        global_tmr_voter(2)(271)  <=    (tmr_registers(0)(271) and tmr_registers(1)(271)) or                                            
                            (tmr_registers(1)(271) and tmr_registers(2)(271)) or                                                       
                            (tmr_registers(0)(271) and tmr_registers(2)(271));                                                         
                                                                                                                                     
        global_tmr_voter(2)(272)  <=    (tmr_registers(0)(272) and tmr_registers(1)(272)) or                                            
                            (tmr_registers(1)(272) and tmr_registers(2)(272)) or                                                       
                            (tmr_registers(0)(272) and tmr_registers(2)(272));                                                         
                                                                                                                                     
        global_tmr_voter(2)(273)  <=    (tmr_registers(0)(273) and tmr_registers(1)(273)) or                                            
                            (tmr_registers(1)(273) and tmr_registers(2)(273)) or                                                       
                            (tmr_registers(0)(273) and tmr_registers(2)(273));                                                         
                                                                                                                                     
        global_tmr_voter(2)(274)  <=    (tmr_registers(0)(274) and tmr_registers(1)(274)) or                                            
                            (tmr_registers(1)(274) and tmr_registers(2)(274)) or                                                       
                            (tmr_registers(0)(274) and tmr_registers(2)(274));                                                         
                                                                                                                                     
        global_tmr_voter(2)(275)  <=    (tmr_registers(0)(275) and tmr_registers(1)(275)) or                                            
                            (tmr_registers(1)(275) and tmr_registers(2)(275)) or                                                       
                            (tmr_registers(0)(275) and tmr_registers(2)(275));                                                         
                                                                                                                                     
        global_tmr_voter(2)(276)  <=    (tmr_registers(0)(276) and tmr_registers(1)(276)) or                                            
                            (tmr_registers(1)(276) and tmr_registers(2)(276)) or                                                       
                            (tmr_registers(0)(276) and tmr_registers(2)(276));                                                         
                                                                                                                                     
        global_tmr_voter(2)(277)  <=    (tmr_registers(0)(277) and tmr_registers(1)(277)) or                                            
                            (tmr_registers(1)(277) and tmr_registers(2)(277)) or                                                       
                            (tmr_registers(0)(277) and tmr_registers(2)(277));                                                         
                                                                                                                                     
        global_tmr_voter(2)(278)  <=    (tmr_registers(0)(278) and tmr_registers(1)(278)) or                                            
                            (tmr_registers(1)(278) and tmr_registers(2)(278)) or                                                       
                            (tmr_registers(0)(278) and tmr_registers(2)(278));                                                         
                                                                                                                                     
        global_tmr_voter(2)(279)  <=    (tmr_registers(0)(279) and tmr_registers(1)(279)) or                                            
                            (tmr_registers(1)(279) and tmr_registers(2)(279)) or                                                       
                            (tmr_registers(0)(279) and tmr_registers(2)(279));                                                         
                                                                                                                                     
        global_tmr_voter(2)(280)  <=    (tmr_registers(0)(280) and tmr_registers(1)(280)) or                                            
                            (tmr_registers(1)(280) and tmr_registers(2)(280)) or                                                       
                            (tmr_registers(0)(280) and tmr_registers(2)(280));                                                         
                                                                                                                                     
        global_tmr_voter(2)(281)  <=    (tmr_registers(0)(281) and tmr_registers(1)(281)) or                                            
                            (tmr_registers(1)(281) and tmr_registers(2)(281)) or                                                       
                            (tmr_registers(0)(281) and tmr_registers(2)(281));                                                         
                                                                                                                                     
        global_tmr_voter(2)(282)  <=    (tmr_registers(0)(282) and tmr_registers(1)(282)) or                                            
                            (tmr_registers(1)(282) and tmr_registers(2)(282)) or                                                       
                            (tmr_registers(0)(282) and tmr_registers(2)(282));                                                         
                                                                                                                                     
        global_tmr_voter(2)(283)  <=    (tmr_registers(0)(283) and tmr_registers(1)(283)) or                                            
                            (tmr_registers(1)(283) and tmr_registers(2)(283)) or                                                       
                            (tmr_registers(0)(283) and tmr_registers(2)(283));                                                         
                                                                                                                                     
        global_tmr_voter(2)(284)  <=    (tmr_registers(0)(284) and tmr_registers(1)(284)) or                                            
                            (tmr_registers(1)(284) and tmr_registers(2)(284)) or                                                       
                            (tmr_registers(0)(284) and tmr_registers(2)(284));                                                         
                                                                                                                                     
        global_tmr_voter(2)(285)  <=    (tmr_registers(0)(285) and tmr_registers(1)(285)) or                                            
                            (tmr_registers(1)(285) and tmr_registers(2)(285)) or                                                       
                            (tmr_registers(0)(285) and tmr_registers(2)(285));                                                         
                                                                                                                                     
        global_tmr_voter(2)(286)  <=    (tmr_registers(0)(286) and tmr_registers(1)(286)) or                                            
                            (tmr_registers(1)(286) and tmr_registers(2)(286)) or                                                       
                            (tmr_registers(0)(286) and tmr_registers(2)(286));                                                         
                                                                                                                                     
        global_tmr_voter(2)(287)  <=    (tmr_registers(0)(287) and tmr_registers(1)(287)) or                                            
                            (tmr_registers(1)(287) and tmr_registers(2)(287)) or                                                       
                            (tmr_registers(0)(287) and tmr_registers(2)(287));                                                         
                                                                                                                                     
        global_tmr_voter(2)(288)  <=    (tmr_registers(0)(288) and tmr_registers(1)(288)) or                                            
                            (tmr_registers(1)(288) and tmr_registers(2)(288)) or                                                       
                            (tmr_registers(0)(288) and tmr_registers(2)(288));                                                         
                                                                                                                                     
        global_tmr_voter(2)(289)  <=    (tmr_registers(0)(289) and tmr_registers(1)(289)) or                                            
                            (tmr_registers(1)(289) and tmr_registers(2)(289)) or                                                       
                            (tmr_registers(0)(289) and tmr_registers(2)(289));                                                         
                                                                                                                                     
        global_tmr_voter(2)(290)  <=    (tmr_registers(0)(290) and tmr_registers(1)(290)) or                                            
                            (tmr_registers(1)(290) and tmr_registers(2)(290)) or                                                       
                            (tmr_registers(0)(290) and tmr_registers(2)(290));                                                         
                                                                                                                                     
        global_tmr_voter(2)(291)  <=    (tmr_registers(0)(291) and tmr_registers(1)(291)) or                                            
                            (tmr_registers(1)(291) and tmr_registers(2)(291)) or                                                       
                            (tmr_registers(0)(291) and tmr_registers(2)(291));                                                         
                                                                                                                                     
        global_tmr_voter(2)(292)  <=    (tmr_registers(0)(292) and tmr_registers(1)(292)) or                                            
                            (tmr_registers(1)(292) and tmr_registers(2)(292)) or                                                       
                            (tmr_registers(0)(292) and tmr_registers(2)(292));                                                         
                                                                                                                                     
        global_tmr_voter(2)(293)  <=    (tmr_registers(0)(293) and tmr_registers(1)(293)) or                                            
                            (tmr_registers(1)(293) and tmr_registers(2)(293)) or                                                       
                            (tmr_registers(0)(293) and tmr_registers(2)(293));                                                         
                                                                                                                                     
        global_tmr_voter(2)(294)  <=    (tmr_registers(0)(294) and tmr_registers(1)(294)) or                                            
                            (tmr_registers(1)(294) and tmr_registers(2)(294)) or                                                       
                            (tmr_registers(0)(294) and tmr_registers(2)(294));                                                         
                                                                                                                                     
        global_tmr_voter(2)(295)  <=    (tmr_registers(0)(295) and tmr_registers(1)(295)) or                                            
                            (tmr_registers(1)(295) and tmr_registers(2)(295)) or                                                       
                            (tmr_registers(0)(295) and tmr_registers(2)(295));                                                         
                                                                                                                                     
        global_tmr_voter(2)(296)  <=    (tmr_registers(0)(296) and tmr_registers(1)(296)) or                                            
                            (tmr_registers(1)(296) and tmr_registers(2)(296)) or                                                       
                            (tmr_registers(0)(296) and tmr_registers(2)(296));                                                         
                                                                                                                                     
        global_tmr_voter(2)(297)  <=    (tmr_registers(0)(297) and tmr_registers(1)(297)) or                                            
                            (tmr_registers(1)(297) and tmr_registers(2)(297)) or                                                       
                            (tmr_registers(0)(297) and tmr_registers(2)(297));                                                         
                                                                                                                                     
        global_tmr_voter(2)(298)  <=    (tmr_registers(0)(298) and tmr_registers(1)(298)) or                                            
                            (tmr_registers(1)(298) and tmr_registers(2)(298)) or                                                       
                            (tmr_registers(0)(298) and tmr_registers(2)(298));                                                         
                                                                                                                                     
        global_tmr_voter(2)(299)  <=    (tmr_registers(0)(299) and tmr_registers(1)(299)) or                                            
                            (tmr_registers(1)(299) and tmr_registers(2)(299)) or                                                       
                            (tmr_registers(0)(299) and tmr_registers(2)(299));                                                         
                                                                                                                                     
        global_tmr_voter(2)(300)  <=    (tmr_registers(0)(300) and tmr_registers(1)(300)) or                                            
                            (tmr_registers(1)(300) and tmr_registers(2)(300)) or                                                       
                            (tmr_registers(0)(300) and tmr_registers(2)(300));                                                         
                                                                                                                                     
        global_tmr_voter(2)(301)  <=    (tmr_registers(0)(301) and tmr_registers(1)(301)) or                                            
                            (tmr_registers(1)(301) and tmr_registers(2)(301)) or                                                       
                            (tmr_registers(0)(301) and tmr_registers(2)(301));                                                         
                                                                                                                                     
        global_tmr_voter(2)(302)  <=    (tmr_registers(0)(302) and tmr_registers(1)(302)) or                                            
                            (tmr_registers(1)(302) and tmr_registers(2)(302)) or                                                       
                            (tmr_registers(0)(302) and tmr_registers(2)(302));                                                         
                                                                                                                                     
        global_tmr_voter(2)(303)  <=    (tmr_registers(0)(303) and tmr_registers(1)(303)) or                                            
                            (tmr_registers(1)(303) and tmr_registers(2)(303)) or                                                       
                            (tmr_registers(0)(303) and tmr_registers(2)(303));                                                         
                                                                                                                                     
        global_tmr_voter(2)(304)  <=    (tmr_registers(0)(304) and tmr_registers(1)(304)) or                                            
                            (tmr_registers(1)(304) and tmr_registers(2)(304)) or                                                       
                            (tmr_registers(0)(304) and tmr_registers(2)(304));                                                         
                                                                                                                                     
        global_tmr_voter(2)(305)  <=    (tmr_registers(0)(305) and tmr_registers(1)(305)) or                                            
                            (tmr_registers(1)(305) and tmr_registers(2)(305)) or                                                       
                            (tmr_registers(0)(305) and tmr_registers(2)(305));                                                         
                                                                                                                                     
        global_tmr_voter(2)(306)  <=    (tmr_registers(0)(306) and tmr_registers(1)(306)) or                                            
                            (tmr_registers(1)(306) and tmr_registers(2)(306)) or                                                       
                            (tmr_registers(0)(306) and tmr_registers(2)(306));                                                         
                                                                                                                                     
        global_tmr_voter(2)(307)  <=    (tmr_registers(0)(307) and tmr_registers(1)(307)) or                                            
                            (tmr_registers(1)(307) and tmr_registers(2)(307)) or                                                       
                            (tmr_registers(0)(307) and tmr_registers(2)(307));                                                         
                                                                                                                                     
        global_tmr_voter(2)(308)  <=    (tmr_registers(0)(308) and tmr_registers(1)(308)) or                                            
                            (tmr_registers(1)(308) and tmr_registers(2)(308)) or                                                       
                            (tmr_registers(0)(308) and tmr_registers(2)(308));                                                         
                                                                                                                                     
        global_tmr_voter(2)(309)  <=    (tmr_registers(0)(309) and tmr_registers(1)(309)) or                                            
                            (tmr_registers(1)(309) and tmr_registers(2)(309)) or                                                       
                            (tmr_registers(0)(309) and tmr_registers(2)(309));                                                         
                                                                                                                                     
        global_tmr_voter(2)(310)  <=    (tmr_registers(0)(310) and tmr_registers(1)(310)) or                                            
                            (tmr_registers(1)(310) and tmr_registers(2)(310)) or                                                       
                            (tmr_registers(0)(310) and tmr_registers(2)(310));                                                         
                                                                                                                                     
        global_tmr_voter(2)(311)  <=    (tmr_registers(0)(311) and tmr_registers(1)(311)) or                                            
                            (tmr_registers(1)(311) and tmr_registers(2)(311)) or                                                       
                            (tmr_registers(0)(311) and tmr_registers(2)(311));                                                         
                                                                                                                                     
        global_tmr_voter(2)(312)  <=    (tmr_registers(0)(312) and tmr_registers(1)(312)) or                                            
                            (tmr_registers(1)(312) and tmr_registers(2)(312)) or                                                       
                            (tmr_registers(0)(312) and tmr_registers(2)(312));                                                         
                                                                                                                                     
        global_tmr_voter(2)(313)  <=    (tmr_registers(0)(313) and tmr_registers(1)(313)) or                                            
                            (tmr_registers(1)(313) and tmr_registers(2)(313)) or                                                       
                            (tmr_registers(0)(313) and tmr_registers(2)(313));                                                         
                                                                                                                                     
        global_tmr_voter(2)(314)  <=    (tmr_registers(0)(314) and tmr_registers(1)(314)) or                                            
                            (tmr_registers(1)(314) and tmr_registers(2)(314)) or                                                       
                            (tmr_registers(0)(314) and tmr_registers(2)(314));                                                         
                                                                                                                                     
        global_tmr_voter(2)(315)  <=    (tmr_registers(0)(315) and tmr_registers(1)(315)) or                                            
                            (tmr_registers(1)(315) and tmr_registers(2)(315)) or                                                       
                            (tmr_registers(0)(315) and tmr_registers(2)(315));                                                         
                                                                                                                                     
        global_tmr_voter(2)(316)  <=    (tmr_registers(0)(316) and tmr_registers(1)(316)) or                                            
                            (tmr_registers(1)(316) and tmr_registers(2)(316)) or                                                       
                            (tmr_registers(0)(316) and tmr_registers(2)(316));                                                         
                                                                                                                                     
        global_tmr_voter(2)(317)  <=    (tmr_registers(0)(317) and tmr_registers(1)(317)) or                                            
                            (tmr_registers(1)(317) and tmr_registers(2)(317)) or                                                       
                            (tmr_registers(0)(317) and tmr_registers(2)(317));                                                         
                                                                                                                                     
        global_tmr_voter(2)(318)  <=    (tmr_registers(0)(318) and tmr_registers(1)(318)) or                                            
                            (tmr_registers(1)(318) and tmr_registers(2)(318)) or                                                       
                            (tmr_registers(0)(318) and tmr_registers(2)(318));                                                         
                                                                                                                                     
        global_tmr_voter(2)(319)  <=    (tmr_registers(0)(319) and tmr_registers(1)(319)) or                                            
                            (tmr_registers(1)(319) and tmr_registers(2)(319)) or                                                       
                            (tmr_registers(0)(319) and tmr_registers(2)(319));                                                         
                                                                                                                                     
        global_tmr_voter(2)(320)  <=    (tmr_registers(0)(320) and tmr_registers(1)(320)) or                                            
                            (tmr_registers(1)(320) and tmr_registers(2)(320)) or                                                       
                            (tmr_registers(0)(320) and tmr_registers(2)(320));                                                         
                                                                                                                                     
        global_tmr_voter(2)(321)  <=    (tmr_registers(0)(321) and tmr_registers(1)(321)) or                                            
                            (tmr_registers(1)(321) and tmr_registers(2)(321)) or                                                       
                            (tmr_registers(0)(321) and tmr_registers(2)(321));                                                         
                                                                                                                                     
        global_tmr_voter(2)(322)  <=    (tmr_registers(0)(322) and tmr_registers(1)(322)) or                                            
                            (tmr_registers(1)(322) and tmr_registers(2)(322)) or                                                       
                            (tmr_registers(0)(322) and tmr_registers(2)(322));                                                         
                                                                                                                                     
        global_tmr_voter(2)(323)  <=    (tmr_registers(0)(323) and tmr_registers(1)(323)) or                                            
                            (tmr_registers(1)(323) and tmr_registers(2)(323)) or                                                       
                            (tmr_registers(0)(323) and tmr_registers(2)(323));                                                         
                                                                                                                                     
        global_tmr_voter(2)(324)  <=    (tmr_registers(0)(324) and tmr_registers(1)(324)) or                                            
                            (tmr_registers(1)(324) and tmr_registers(2)(324)) or                                                       
                            (tmr_registers(0)(324) and tmr_registers(2)(324));                                                         
                                                                                                                                     
        global_tmr_voter(2)(325)  <=    (tmr_registers(0)(325) and tmr_registers(1)(325)) or                                            
                            (tmr_registers(1)(325) and tmr_registers(2)(325)) or                                                       
                            (tmr_registers(0)(325) and tmr_registers(2)(325));                                                         
                                                                                                                                     
        global_tmr_voter(2)(326)  <=    (tmr_registers(0)(326) and tmr_registers(1)(326)) or                                            
                            (tmr_registers(1)(326) and tmr_registers(2)(326)) or                                                       
                            (tmr_registers(0)(326) and tmr_registers(2)(326));                                                         
                                                                                                                                     
        global_tmr_voter(2)(327)  <=    (tmr_registers(0)(327) and tmr_registers(1)(327)) or                                            
                            (tmr_registers(1)(327) and tmr_registers(2)(327)) or                                                       
                            (tmr_registers(0)(327) and tmr_registers(2)(327));                                                         
                                                                                                                                     
        global_tmr_voter(2)(328)  <=    (tmr_registers(0)(328) and tmr_registers(1)(328)) or                                            
                            (tmr_registers(1)(328) and tmr_registers(2)(328)) or                                                       
                            (tmr_registers(0)(328) and tmr_registers(2)(328));                                                         
                                                                                                                                     
        global_tmr_voter(2)(329)  <=    (tmr_registers(0)(329) and tmr_registers(1)(329)) or                                            
                            (tmr_registers(1)(329) and tmr_registers(2)(329)) or                                                       
                            (tmr_registers(0)(329) and tmr_registers(2)(329));                                                         
                                                                                                                                     
        global_tmr_voter(2)(330)  <=    (tmr_registers(0)(330) and tmr_registers(1)(330)) or                                            
                            (tmr_registers(1)(330) and tmr_registers(2)(330)) or                                                       
                            (tmr_registers(0)(330) and tmr_registers(2)(330));                                                         
                                                                                                                                     
        global_tmr_voter(2)(331)  <=    (tmr_registers(0)(331) and tmr_registers(1)(331)) or                                            
                            (tmr_registers(1)(331) and tmr_registers(2)(331)) or                                                       
                            (tmr_registers(0)(331) and tmr_registers(2)(331));                                                         
                                                                                                                                     
        global_tmr_voter(2)(332)  <=    (tmr_registers(0)(332) and tmr_registers(1)(332)) or                                            
                            (tmr_registers(1)(332) and tmr_registers(2)(332)) or                                                       
                            (tmr_registers(0)(332) and tmr_registers(2)(332));                                                         
                                                                                                                                     
        global_tmr_voter(2)(333)  <=    (tmr_registers(0)(333) and tmr_registers(1)(333)) or                                            
                            (tmr_registers(1)(333) and tmr_registers(2)(333)) or                                                       
                            (tmr_registers(0)(333) and tmr_registers(2)(333));                                                         
                                                                                                                                     
        global_tmr_voter(2)(334)  <=    (tmr_registers(0)(334) and tmr_registers(1)(334)) or                                            
                            (tmr_registers(1)(334) and tmr_registers(2)(334)) or                                                       
                            (tmr_registers(0)(334) and tmr_registers(2)(334));                                                         
                                                                                                                                     
        global_tmr_voter(2)(335)  <=    (tmr_registers(0)(335) and tmr_registers(1)(335)) or                                            
                            (tmr_registers(1)(335) and tmr_registers(2)(335)) or                                                       
                            (tmr_registers(0)(335) and tmr_registers(2)(335));                                                         
                                                                                                                                     
        global_tmr_voter(2)(336)  <=    (tmr_registers(0)(336) and tmr_registers(1)(336)) or                                            
                            (tmr_registers(1)(336) and tmr_registers(2)(336)) or                                                       
                            (tmr_registers(0)(336) and tmr_registers(2)(336));                                                         
                                                                                                                                     
        global_tmr_voter(2)(337)  <=    (tmr_registers(0)(337) and tmr_registers(1)(337)) or                                            
                            (tmr_registers(1)(337) and tmr_registers(2)(337)) or                                                       
                            (tmr_registers(0)(337) and tmr_registers(2)(337));                                                         
                                                                                                                                     
        global_tmr_voter(2)(338)  <=    (tmr_registers(0)(338) and tmr_registers(1)(338)) or                                            
                            (tmr_registers(1)(338) and tmr_registers(2)(338)) or                                                       
                            (tmr_registers(0)(338) and tmr_registers(2)(338));                                                         
                                                                                                                                     
        global_tmr_voter(2)(339)  <=    (tmr_registers(0)(339) and tmr_registers(1)(339)) or                                            
                            (tmr_registers(1)(339) and tmr_registers(2)(339)) or                                                       
                            (tmr_registers(0)(339) and tmr_registers(2)(339));                                                         
                                                                                                                                     
        global_tmr_voter(2)(340)  <=    (tmr_registers(0)(340) and tmr_registers(1)(340)) or                                            
                            (tmr_registers(1)(340) and tmr_registers(2)(340)) or                                                       
                            (tmr_registers(0)(340) and tmr_registers(2)(340));                                                         
                                                                                                                                     
        global_tmr_voter(2)(341)  <=    (tmr_registers(0)(341) and tmr_registers(1)(341)) or                                            
                            (tmr_registers(1)(341) and tmr_registers(2)(341)) or                                                       
                            (tmr_registers(0)(341) and tmr_registers(2)(341));                                                         
                                                                                                                                     
        global_tmr_voter(2)(342)  <=    (tmr_registers(0)(342) and tmr_registers(1)(342)) or                                            
                            (tmr_registers(1)(342) and tmr_registers(2)(342)) or                                                       
                            (tmr_registers(0)(342) and tmr_registers(2)(342));                                                         
                                                                                                                                     
        global_tmr_voter(2)(343)  <=    (tmr_registers(0)(343) and tmr_registers(1)(343)) or                                            
                            (tmr_registers(1)(343) and tmr_registers(2)(343)) or                                                       
                            (tmr_registers(0)(343) and tmr_registers(2)(343));                                                         
                                                                                                                                     
        global_tmr_voter(2)(344)  <=    (tmr_registers(0)(344) and tmr_registers(1)(344)) or                                            
                            (tmr_registers(1)(344) and tmr_registers(2)(344)) or                                                       
                            (tmr_registers(0)(344) and tmr_registers(2)(344));                                                         
                                                                                                                                     
        global_tmr_voter(2)(345)  <=    (tmr_registers(0)(345) and tmr_registers(1)(345)) or                                            
                            (tmr_registers(1)(345) and tmr_registers(2)(345)) or                                                       
                            (tmr_registers(0)(345) and tmr_registers(2)(345));                                                         
                                                                                                                                     
        global_tmr_voter(2)(346)  <=    (tmr_registers(0)(346) and tmr_registers(1)(346)) or                                            
                            (tmr_registers(1)(346) and tmr_registers(2)(346)) or                                                       
                            (tmr_registers(0)(346) and tmr_registers(2)(346));                                                         
                                                                                                                                     
        global_tmr_voter(2)(347)  <=    (tmr_registers(0)(347) and tmr_registers(1)(347)) or                                            
                            (tmr_registers(1)(347) and tmr_registers(2)(347)) or                                                       
                            (tmr_registers(0)(347) and tmr_registers(2)(347));                                                         
                                                                                                                                     
        global_tmr_voter(2)(348)  <=    (tmr_registers(0)(348) and tmr_registers(1)(348)) or                                            
                            (tmr_registers(1)(348) and tmr_registers(2)(348)) or                                                       
                            (tmr_registers(0)(348) and tmr_registers(2)(348));                                                         
                                                                                                                                     
        global_tmr_voter(2)(349)  <=    (tmr_registers(0)(349) and tmr_registers(1)(349)) or                                            
                            (tmr_registers(1)(349) and tmr_registers(2)(349)) or                                                       
                            (tmr_registers(0)(349) and tmr_registers(2)(349));                                                         
                                                                                                                                     
        global_tmr_voter(2)(350)  <=    (tmr_registers(0)(350) and tmr_registers(1)(350)) or                                            
                            (tmr_registers(1)(350) and tmr_registers(2)(350)) or                                                       
                            (tmr_registers(0)(350) and tmr_registers(2)(350));                                                         
                                                                                                                                     
        global_tmr_voter(2)(351)  <=    (tmr_registers(0)(351) and tmr_registers(1)(351)) or                                            
                            (tmr_registers(1)(351) and tmr_registers(2)(351)) or                                                       
                            (tmr_registers(0)(351) and tmr_registers(2)(351));                                                         
                                                                                                                                     
        global_tmr_voter(2)(352)  <=    (tmr_registers(0)(352) and tmr_registers(1)(352)) or                                            
                            (tmr_registers(1)(352) and tmr_registers(2)(352)) or                                                       
                            (tmr_registers(0)(352) and tmr_registers(2)(352));                                                         
                                                                                                                                     
        global_tmr_voter(2)(353)  <=    (tmr_registers(0)(353) and tmr_registers(1)(353)) or                                            
                            (tmr_registers(1)(353) and tmr_registers(2)(353)) or                                                       
                            (tmr_registers(0)(353) and tmr_registers(2)(353));                                                         
                                                                                                                                     
        global_tmr_voter(2)(354)  <=    (tmr_registers(0)(354) and tmr_registers(1)(354)) or                                            
                            (tmr_registers(1)(354) and tmr_registers(2)(354)) or                                                       
                            (tmr_registers(0)(354) and tmr_registers(2)(354));                                                         
                                                                                                                                     
        global_tmr_voter(2)(355)  <=    (tmr_registers(0)(355) and tmr_registers(1)(355)) or                                            
                            (tmr_registers(1)(355) and tmr_registers(2)(355)) or                                                       
                            (tmr_registers(0)(355) and tmr_registers(2)(355));                                                         
                                                                                                                                     
        global_tmr_voter(2)(356)  <=    (tmr_registers(0)(356) and tmr_registers(1)(356)) or                                            
                            (tmr_registers(1)(356) and tmr_registers(2)(356)) or                                                       
                            (tmr_registers(0)(356) and tmr_registers(2)(356));                                                         
                                                                                                                                     
        global_tmr_voter(2)(357)  <=    (tmr_registers(0)(357) and tmr_registers(1)(357)) or                                            
                            (tmr_registers(1)(357) and tmr_registers(2)(357)) or                                                       
                            (tmr_registers(0)(357) and tmr_registers(2)(357));                                                         
                                                                                                                                     
        global_tmr_voter(2)(358)  <=    (tmr_registers(0)(358) and tmr_registers(1)(358)) or                                            
                            (tmr_registers(1)(358) and tmr_registers(2)(358)) or                                                       
                            (tmr_registers(0)(358) and tmr_registers(2)(358));                                                         
                                                                                                                                     
        global_tmr_voter(2)(359)  <=    (tmr_registers(0)(359) and tmr_registers(1)(359)) or                                            
                            (tmr_registers(1)(359) and tmr_registers(2)(359)) or                                                       
                            (tmr_registers(0)(359) and tmr_registers(2)(359));                                                         
                                                                                                                                     
        global_tmr_voter(2)(360)  <=    (tmr_registers(0)(360) and tmr_registers(1)(360)) or                                            
                            (tmr_registers(1)(360) and tmr_registers(2)(360)) or                                                       
                            (tmr_registers(0)(360) and tmr_registers(2)(360));                                                         
                                                                                                                                     
        global_tmr_voter(2)(361)  <=    (tmr_registers(0)(361) and tmr_registers(1)(361)) or                                            
                            (tmr_registers(1)(361) and tmr_registers(2)(361)) or                                                       
                            (tmr_registers(0)(361) and tmr_registers(2)(361));                                                         
                                                                                                                                     
        global_tmr_voter(2)(362)  <=    (tmr_registers(0)(362) and tmr_registers(1)(362)) or                                            
                            (tmr_registers(1)(362) and tmr_registers(2)(362)) or                                                       
                            (tmr_registers(0)(362) and tmr_registers(2)(362));                                                         
                                                                                                                                     
        global_tmr_voter(2)(363)  <=    (tmr_registers(0)(363) and tmr_registers(1)(363)) or                                            
                            (tmr_registers(1)(363) and tmr_registers(2)(363)) or                                                       
                            (tmr_registers(0)(363) and tmr_registers(2)(363));                                                         
                                                                                                                                     
        global_tmr_voter(2)(364)  <=    (tmr_registers(0)(364) and tmr_registers(1)(364)) or                                            
                            (tmr_registers(1)(364) and tmr_registers(2)(364)) or                                                       
                            (tmr_registers(0)(364) and tmr_registers(2)(364));                                                         
                                                                                                                                     
        global_tmr_voter(2)(365)  <=    (tmr_registers(0)(365) and tmr_registers(1)(365)) or                                            
                            (tmr_registers(1)(365) and tmr_registers(2)(365)) or                                                       
                            (tmr_registers(0)(365) and tmr_registers(2)(365));                                                         
                                                                                                                                     
        global_tmr_voter(2)(366)  <=    (tmr_registers(0)(366) and tmr_registers(1)(366)) or                                            
                            (tmr_registers(1)(366) and tmr_registers(2)(366)) or                                                       
                            (tmr_registers(0)(366) and tmr_registers(2)(366));                                                         
                                                                                                                                     
        global_tmr_voter(2)(367)  <=    (tmr_registers(0)(367) and tmr_registers(1)(367)) or                                            
                            (tmr_registers(1)(367) and tmr_registers(2)(367)) or                                                       
                            (tmr_registers(0)(367) and tmr_registers(2)(367));                                                         
                                                                                                                                     
        global_tmr_voter(2)(368)  <=    (tmr_registers(0)(368) and tmr_registers(1)(368)) or                                            
                            (tmr_registers(1)(368) and tmr_registers(2)(368)) or                                                       
                            (tmr_registers(0)(368) and tmr_registers(2)(368));                                                         
                                                                                                                                     
        global_tmr_voter(2)(369)  <=    (tmr_registers(0)(369) and tmr_registers(1)(369)) or                                            
                            (tmr_registers(1)(369) and tmr_registers(2)(369)) or                                                       
                            (tmr_registers(0)(369) and tmr_registers(2)(369));                                                         
                                                                                                                                     
        global_tmr_voter(2)(370)  <=    (tmr_registers(0)(370) and tmr_registers(1)(370)) or                                            
                            (tmr_registers(1)(370) and tmr_registers(2)(370)) or                                                       
                            (tmr_registers(0)(370) and tmr_registers(2)(370));                                                         
                                                                                                                                     
        global_tmr_voter(2)(371)  <=    (tmr_registers(0)(371) and tmr_registers(1)(371)) or                                            
                            (tmr_registers(1)(371) and tmr_registers(2)(371)) or                                                       
                            (tmr_registers(0)(371) and tmr_registers(2)(371));                                                         
                                                                                                                                     
        global_tmr_voter(2)(372)  <=    (tmr_registers(0)(372) and tmr_registers(1)(372)) or                                            
                            (tmr_registers(1)(372) and tmr_registers(2)(372)) or                                                       
                            (tmr_registers(0)(372) and tmr_registers(2)(372));                                                         
                                                                                                                                     
        global_tmr_voter(2)(373)  <=    (tmr_registers(0)(373) and tmr_registers(1)(373)) or                                            
                            (tmr_registers(1)(373) and tmr_registers(2)(373)) or                                                       
                            (tmr_registers(0)(373) and tmr_registers(2)(373));                                                         
                                                                                                                                     
        global_tmr_voter(2)(374)  <=    (tmr_registers(0)(374) and tmr_registers(1)(374)) or                                            
                            (tmr_registers(1)(374) and tmr_registers(2)(374)) or                                                       
                            (tmr_registers(0)(374) and tmr_registers(2)(374));                                                         
                                                                                                                                     
        global_tmr_voter(2)(375)  <=    (tmr_registers(0)(375) and tmr_registers(1)(375)) or                                            
                            (tmr_registers(1)(375) and tmr_registers(2)(375)) or                                                       
                            (tmr_registers(0)(375) and tmr_registers(2)(375));                                                         
                                                                                                                                     
        global_tmr_voter(2)(376)  <=    (tmr_registers(0)(376) and tmr_registers(1)(376)) or                                            
                            (tmr_registers(1)(376) and tmr_registers(2)(376)) or                                                       
                            (tmr_registers(0)(376) and tmr_registers(2)(376));                                                         
                                                                                                                                     
        global_tmr_voter(2)(377)  <=    (tmr_registers(0)(377) and tmr_registers(1)(377)) or                                            
                            (tmr_registers(1)(377) and tmr_registers(2)(377)) or                                                       
                            (tmr_registers(0)(377) and tmr_registers(2)(377));                                                         
                                                                                                                                     
        global_tmr_voter(2)(378)  <=    (tmr_registers(0)(378) and tmr_registers(1)(378)) or                                            
                            (tmr_registers(1)(378) and tmr_registers(2)(378)) or                                                       
                            (tmr_registers(0)(378) and tmr_registers(2)(378));                                                         
                                                                                                                                     
        global_tmr_voter(2)(379)  <=    (tmr_registers(0)(379) and tmr_registers(1)(379)) or                                            
                            (tmr_registers(1)(379) and tmr_registers(2)(379)) or                                                       
                            (tmr_registers(0)(379) and tmr_registers(2)(379));                                                         
                                                                                                                                     
        global_tmr_voter(2)(380)  <=    (tmr_registers(0)(380) and tmr_registers(1)(380)) or                                            
                            (tmr_registers(1)(380) and tmr_registers(2)(380)) or                                                       
                            (tmr_registers(0)(380) and tmr_registers(2)(380));                                                         
                                                                                                                                     
        global_tmr_voter(2)(381)  <=    (tmr_registers(0)(381) and tmr_registers(1)(381)) or                                            
                            (tmr_registers(1)(381) and tmr_registers(2)(381)) or                                                       
                            (tmr_registers(0)(381) and tmr_registers(2)(381));                                                         
                                                                                                                                     
        global_tmr_voter(2)(382)  <=    (tmr_registers(0)(382) and tmr_registers(1)(382)) or                                            
                            (tmr_registers(1)(382) and tmr_registers(2)(382)) or                                                       
                            (tmr_registers(0)(382) and tmr_registers(2)(382));                                                         
                                                                                                                                     
        global_tmr_voter(2)(383)  <=    (tmr_registers(0)(383) and tmr_registers(1)(383)) or                                            
                            (tmr_registers(1)(383) and tmr_registers(2)(383)) or                                                       
                            (tmr_registers(0)(383) and tmr_registers(2)(383));                                                         
                                                                                                                                     
        global_tmr_voter(2)(384)  <=    (tmr_registers(0)(384) and tmr_registers(1)(384)) or                                            
                            (tmr_registers(1)(384) and tmr_registers(2)(384)) or                                                       
                            (tmr_registers(0)(384) and tmr_registers(2)(384));                                                         
                                                                                                                                     
        global_tmr_voter(2)(385)  <=    (tmr_registers(0)(385) and tmr_registers(1)(385)) or                                            
                            (tmr_registers(1)(385) and tmr_registers(2)(385)) or                                                       
                            (tmr_registers(0)(385) and tmr_registers(2)(385));                                                         
                                                                                                                                     
        global_tmr_voter(2)(386)  <=    (tmr_registers(0)(386) and tmr_registers(1)(386)) or                                            
                            (tmr_registers(1)(386) and tmr_registers(2)(386)) or                                                       
                            (tmr_registers(0)(386) and tmr_registers(2)(386));                                                         
                                                                                                                                     
        global_tmr_voter(2)(387)  <=    (tmr_registers(0)(387) and tmr_registers(1)(387)) or                                            
                            (tmr_registers(1)(387) and tmr_registers(2)(387)) or                                                       
                            (tmr_registers(0)(387) and tmr_registers(2)(387));                                                         
                                                                                                                                     
        global_tmr_voter(2)(388)  <=    (tmr_registers(0)(388) and tmr_registers(1)(388)) or                                            
                            (tmr_registers(1)(388) and tmr_registers(2)(388)) or                                                       
                            (tmr_registers(0)(388) and tmr_registers(2)(388));                                                         
                                                                                                                                     
        global_tmr_voter(2)(389)  <=    (tmr_registers(0)(389) and tmr_registers(1)(389)) or                                            
                            (tmr_registers(1)(389) and tmr_registers(2)(389)) or                                                       
                            (tmr_registers(0)(389) and tmr_registers(2)(389));                                                         
                                                                                                                                     
        global_tmr_voter(2)(390)  <=    (tmr_registers(0)(390) and tmr_registers(1)(390)) or                                            
                            (tmr_registers(1)(390) and tmr_registers(2)(390)) or                                                       
                            (tmr_registers(0)(390) and tmr_registers(2)(390));                                                         
                                                                                                                                     
        global_tmr_voter(2)(391)  <=    (tmr_registers(0)(391) and tmr_registers(1)(391)) or                                            
                            (tmr_registers(1)(391) and tmr_registers(2)(391)) or                                                       
                            (tmr_registers(0)(391) and tmr_registers(2)(391));                                                         
                                                                                                                                     
        global_tmr_voter(2)(392)  <=    (tmr_registers(0)(392) and tmr_registers(1)(392)) or                                            
                            (tmr_registers(1)(392) and tmr_registers(2)(392)) or                                                       
                            (tmr_registers(0)(392) and tmr_registers(2)(392));                                                         
                                                                                                                                     
        global_tmr_voter(2)(393)  <=    (tmr_registers(0)(393) and tmr_registers(1)(393)) or                                            
                            (tmr_registers(1)(393) and tmr_registers(2)(393)) or                                                       
                            (tmr_registers(0)(393) and tmr_registers(2)(393));                                                         
                                                                                                                                     
        global_tmr_voter(2)(394)  <=    (tmr_registers(0)(394) and tmr_registers(1)(394)) or                                            
                            (tmr_registers(1)(394) and tmr_registers(2)(394)) or                                                       
                            (tmr_registers(0)(394) and tmr_registers(2)(394));                                                         
                                                                                                                                     
        global_tmr_voter(2)(395)  <=    (tmr_registers(0)(395) and tmr_registers(1)(395)) or                                            
                            (tmr_registers(1)(395) and tmr_registers(2)(395)) or                                                       
                            (tmr_registers(0)(395) and tmr_registers(2)(395));                                                         
                                                                                                                                     
        global_tmr_voter(2)(396)  <=    (tmr_registers(0)(396) and tmr_registers(1)(396)) or                                            
                            (tmr_registers(1)(396) and tmr_registers(2)(396)) or                                                       
                            (tmr_registers(0)(396) and tmr_registers(2)(396));                                                         
                                                                                                                                     
        global_tmr_voter(2)(397)  <=    (tmr_registers(0)(397) and tmr_registers(1)(397)) or                                            
                            (tmr_registers(1)(397) and tmr_registers(2)(397)) or                                                       
                            (tmr_registers(0)(397) and tmr_registers(2)(397));                                                         
                                                                                                                                     
        global_tmr_voter(2)(398)  <=    (tmr_registers(0)(398) and tmr_registers(1)(398)) or                                            
                            (tmr_registers(1)(398) and tmr_registers(2)(398)) or                                                       
                            (tmr_registers(0)(398) and tmr_registers(2)(398));                                                         
                                                                                                                                     
        global_tmr_voter(2)(399)  <=    (tmr_registers(0)(399) and tmr_registers(1)(399)) or                                            
                            (tmr_registers(1)(399) and tmr_registers(2)(399)) or                                                       
                            (tmr_registers(0)(399) and tmr_registers(2)(399));                                                         
                                                                                                                                     
        global_tmr_voter(2)(400)  <=    (tmr_registers(0)(400) and tmr_registers(1)(400)) or                                            
                            (tmr_registers(1)(400) and tmr_registers(2)(400)) or                                                       
                            (tmr_registers(0)(400) and tmr_registers(2)(400));                                                         
                                                                                                                                     
        global_tmr_voter(2)(401)  <=    (tmr_registers(0)(401) and tmr_registers(1)(401)) or                                            
                            (tmr_registers(1)(401) and tmr_registers(2)(401)) or                                                       
                            (tmr_registers(0)(401) and tmr_registers(2)(401));                                                         
                                                                                                                                     
        global_tmr_voter(2)(402)  <=    (tmr_registers(0)(402) and tmr_registers(1)(402)) or                                            
                            (tmr_registers(1)(402) and tmr_registers(2)(402)) or                                                       
                            (tmr_registers(0)(402) and tmr_registers(2)(402));                                                         
                                                                                                                                     
        global_tmr_voter(2)(403)  <=    (tmr_registers(0)(403) and tmr_registers(1)(403)) or                                            
                            (tmr_registers(1)(403) and tmr_registers(2)(403)) or                                                       
                            (tmr_registers(0)(403) and tmr_registers(2)(403));                                                         
                                                                                                                                     
        global_tmr_voter(2)(404)  <=    (tmr_registers(0)(404) and tmr_registers(1)(404)) or                                            
                            (tmr_registers(1)(404) and tmr_registers(2)(404)) or                                                       
                            (tmr_registers(0)(404) and tmr_registers(2)(404));                                                         
                                                                                                                                     
        global_tmr_voter(2)(405)  <=    (tmr_registers(0)(405) and tmr_registers(1)(405)) or                                            
                            (tmr_registers(1)(405) and tmr_registers(2)(405)) or                                                       
                            (tmr_registers(0)(405) and tmr_registers(2)(405));                                                         
                                                                                                                                     
        global_tmr_voter(2)(406)  <=    (tmr_registers(0)(406) and tmr_registers(1)(406)) or                                            
                            (tmr_registers(1)(406) and tmr_registers(2)(406)) or                                                       
                            (tmr_registers(0)(406) and tmr_registers(2)(406));                                                         
                                                                                                                                     
        global_tmr_voter(2)(407)  <=    (tmr_registers(0)(407) and tmr_registers(1)(407)) or                                            
                            (tmr_registers(1)(407) and tmr_registers(2)(407)) or                                                       
                            (tmr_registers(0)(407) and tmr_registers(2)(407));                                                         
                                                                                                                                     
        global_tmr_voter(2)(408)  <=    (tmr_registers(0)(408) and tmr_registers(1)(408)) or                                            
                            (tmr_registers(1)(408) and tmr_registers(2)(408)) or                                                       
                            (tmr_registers(0)(408) and tmr_registers(2)(408));                                                         
                                                                                                                                     
        global_tmr_voter(2)(409)  <=    (tmr_registers(0)(409) and tmr_registers(1)(409)) or                                            
                            (tmr_registers(1)(409) and tmr_registers(2)(409)) or                                                       
                            (tmr_registers(0)(409) and tmr_registers(2)(409));                                                         
                                                                                                                                     
        global_tmr_voter(2)(410)  <=    (tmr_registers(0)(410) and tmr_registers(1)(410)) or                                            
                            (tmr_registers(1)(410) and tmr_registers(2)(410)) or                                                       
                            (tmr_registers(0)(410) and tmr_registers(2)(410));                                                         
                                                                                                                                     
        global_tmr_voter(2)(411)  <=    (tmr_registers(0)(411) and tmr_registers(1)(411)) or                                            
                            (tmr_registers(1)(411) and tmr_registers(2)(411)) or                                                       
                            (tmr_registers(0)(411) and tmr_registers(2)(411));                                                         
                                                                                                                                     
        global_tmr_voter(2)(412)  <=    (tmr_registers(0)(412) and tmr_registers(1)(412)) or                                            
                            (tmr_registers(1)(412) and tmr_registers(2)(412)) or                                                       
                            (tmr_registers(0)(412) and tmr_registers(2)(412));                                                         
                                                                                                                                     
        global_tmr_voter(2)(413)  <=    (tmr_registers(0)(413) and tmr_registers(1)(413)) or                                            
                            (tmr_registers(1)(413) and tmr_registers(2)(413)) or                                                       
                            (tmr_registers(0)(413) and tmr_registers(2)(413));                                                         
                                                                                                                                     
        global_tmr_voter(2)(414)  <=    (tmr_registers(0)(414) and tmr_registers(1)(414)) or                                            
                            (tmr_registers(1)(414) and tmr_registers(2)(414)) or                                                       
                            (tmr_registers(0)(414) and tmr_registers(2)(414));                                                         
                                                                                                                                     
        global_tmr_voter(2)(415)  <=    (tmr_registers(0)(415) and tmr_registers(1)(415)) or                                            
                            (tmr_registers(1)(415) and tmr_registers(2)(415)) or                                                       
                            (tmr_registers(0)(415) and tmr_registers(2)(415));                                                         
                                                                                                                                     
        global_tmr_voter(2)(416)  <=    (tmr_registers(0)(416) and tmr_registers(1)(416)) or                                            
                            (tmr_registers(1)(416) and tmr_registers(2)(416)) or                                                       
                            (tmr_registers(0)(416) and tmr_registers(2)(416));                                                         
                                                                                                                                     
        global_tmr_voter(2)(417)  <=    (tmr_registers(0)(417) and tmr_registers(1)(417)) or                                            
                            (tmr_registers(1)(417) and tmr_registers(2)(417)) or                                                       
                            (tmr_registers(0)(417) and tmr_registers(2)(417));                                                         
                                                                                                                                     
        global_tmr_voter(2)(418)  <=    (tmr_registers(0)(418) and tmr_registers(1)(418)) or                                            
                            (tmr_registers(1)(418) and tmr_registers(2)(418)) or                                                       
                            (tmr_registers(0)(418) and tmr_registers(2)(418));                                                         
                                                                                                                                     
        global_tmr_voter(2)(419)  <=    (tmr_registers(0)(419) and tmr_registers(1)(419)) or                                            
                            (tmr_registers(1)(419) and tmr_registers(2)(419)) or                                                       
                            (tmr_registers(0)(419) and tmr_registers(2)(419));                                                         
                                                                                                                                     
        global_tmr_voter(2)(420)  <=    (tmr_registers(0)(420) and tmr_registers(1)(420)) or                                            
                            (tmr_registers(1)(420) and tmr_registers(2)(420)) or                                                       
                            (tmr_registers(0)(420) and tmr_registers(2)(420));                                                         
                                                                                                                                     
        global_tmr_voter(2)(421)  <=    (tmr_registers(0)(421) and tmr_registers(1)(421)) or                                            
                            (tmr_registers(1)(421) and tmr_registers(2)(421)) or                                                       
                            (tmr_registers(0)(421) and tmr_registers(2)(421));                                                         
                                                                                                                                     
        global_tmr_voter(2)(422)  <=    (tmr_registers(0)(422) and tmr_registers(1)(422)) or                                            
                            (tmr_registers(1)(422) and tmr_registers(2)(422)) or                                                       
                            (tmr_registers(0)(422) and tmr_registers(2)(422));                                                         
                                                                                                                                     
        global_tmr_voter(2)(423)  <=    (tmr_registers(0)(423) and tmr_registers(1)(423)) or                                            
                            (tmr_registers(1)(423) and tmr_registers(2)(423)) or                                                       
                            (tmr_registers(0)(423) and tmr_registers(2)(423));                                                         
                                                                                                                                     
        global_tmr_voter(2)(424)  <=    (tmr_registers(0)(424) and tmr_registers(1)(424)) or                                            
                            (tmr_registers(1)(424) and tmr_registers(2)(424)) or                                                       
                            (tmr_registers(0)(424) and tmr_registers(2)(424));                                                         
                                                                                                                                     
        global_tmr_voter(2)(425)  <=    (tmr_registers(0)(425) and tmr_registers(1)(425)) or                                            
                            (tmr_registers(1)(425) and tmr_registers(2)(425)) or                                                       
                            (tmr_registers(0)(425) and tmr_registers(2)(425));                                                         
                                                                                                                                     
        global_tmr_voter(2)(426)  <=    (tmr_registers(0)(426) and tmr_registers(1)(426)) or                                            
                            (tmr_registers(1)(426) and tmr_registers(2)(426)) or                                                       
                            (tmr_registers(0)(426) and tmr_registers(2)(426));                                                         
                                                                                                                                     
        global_tmr_voter(2)(427)  <=    (tmr_registers(0)(427) and tmr_registers(1)(427)) or                                            
                            (tmr_registers(1)(427) and tmr_registers(2)(427)) or                                                       
                            (tmr_registers(0)(427) and tmr_registers(2)(427));                                                         
                                                                                                                                     
        global_tmr_voter(2)(428)  <=    (tmr_registers(0)(428) and tmr_registers(1)(428)) or                                            
                            (tmr_registers(1)(428) and tmr_registers(2)(428)) or                                                       
                            (tmr_registers(0)(428) and tmr_registers(2)(428));                                                         
                                                                                                                                     
        global_tmr_voter(2)(429)  <=    (tmr_registers(0)(429) and tmr_registers(1)(429)) or                                            
                            (tmr_registers(1)(429) and tmr_registers(2)(429)) or                                                       
                            (tmr_registers(0)(429) and tmr_registers(2)(429));                                                         
                                                                                                                                     
        global_tmr_voter(2)(430)  <=    (tmr_registers(0)(430) and tmr_registers(1)(430)) or                                            
                            (tmr_registers(1)(430) and tmr_registers(2)(430)) or                                                       
                            (tmr_registers(0)(430) and tmr_registers(2)(430));                                                         
                                                                                                                                     
        global_tmr_voter(2)(431)  <=    (tmr_registers(0)(431) and tmr_registers(1)(431)) or                                            
                            (tmr_registers(1)(431) and tmr_registers(2)(431)) or                                                       
                            (tmr_registers(0)(431) and tmr_registers(2)(431));                                                         
                                                                                                                                     
        global_tmr_voter(2)(432)  <=    (tmr_registers(0)(432) and tmr_registers(1)(432)) or                                            
                            (tmr_registers(1)(432) and tmr_registers(2)(432)) or                                                       
                            (tmr_registers(0)(432) and tmr_registers(2)(432));                                                         
                                                                                                                                     
        global_tmr_voter(2)(433)  <=    (tmr_registers(0)(433) and tmr_registers(1)(433)) or                                            
                            (tmr_registers(1)(433) and tmr_registers(2)(433)) or                                                       
                            (tmr_registers(0)(433) and tmr_registers(2)(433));                                                         
                                                                                                                                     
        global_tmr_voter(2)(434)  <=    (tmr_registers(0)(434) and tmr_registers(1)(434)) or                                            
                            (tmr_registers(1)(434) and tmr_registers(2)(434)) or                                                       
                            (tmr_registers(0)(434) and tmr_registers(2)(434));                                                         
                                                                                                                                     
        global_tmr_voter(2)(435)  <=    (tmr_registers(0)(435) and tmr_registers(1)(435)) or                                            
                            (tmr_registers(1)(435) and tmr_registers(2)(435)) or                                                       
                            (tmr_registers(0)(435) and tmr_registers(2)(435));                                                         
                                                                                                                                     
        global_tmr_voter(2)(436)  <=    (tmr_registers(0)(436) and tmr_registers(1)(436)) or                                            
                            (tmr_registers(1)(436) and tmr_registers(2)(436)) or                                                       
                            (tmr_registers(0)(436) and tmr_registers(2)(436));                                                         
                                                                                                                                     
        global_tmr_voter(2)(437)  <=    (tmr_registers(0)(437) and tmr_registers(1)(437)) or                                            
                            (tmr_registers(1)(437) and tmr_registers(2)(437)) or                                                       
                            (tmr_registers(0)(437) and tmr_registers(2)(437));                                                         
                                                                                                                                     
        global_tmr_voter(2)(438)  <=    (tmr_registers(0)(438) and tmr_registers(1)(438)) or                                            
                            (tmr_registers(1)(438) and tmr_registers(2)(438)) or                                                       
                            (tmr_registers(0)(438) and tmr_registers(2)(438));                                                         
                                                                                                                                     
        global_tmr_voter(2)(439)  <=    (tmr_registers(0)(439) and tmr_registers(1)(439)) or                                            
                            (tmr_registers(1)(439) and tmr_registers(2)(439)) or                                                       
                            (tmr_registers(0)(439) and tmr_registers(2)(439));                                                         
                                                                                                                                     
        global_tmr_voter(2)(440)  <=    (tmr_registers(0)(440) and tmr_registers(1)(440)) or                                            
                            (tmr_registers(1)(440) and tmr_registers(2)(440)) or                                                       
                            (tmr_registers(0)(440) and tmr_registers(2)(440));                                                         
                                                                                                                                     
        global_tmr_voter(2)(441)  <=    (tmr_registers(0)(441) and tmr_registers(1)(441)) or                                            
                            (tmr_registers(1)(441) and tmr_registers(2)(441)) or                                                       
                            (tmr_registers(0)(441) and tmr_registers(2)(441));                                                         
                                                                                                                                     
        global_tmr_voter(2)(442)  <=    (tmr_registers(0)(442) and tmr_registers(1)(442)) or                                            
                            (tmr_registers(1)(442) and tmr_registers(2)(442)) or                                                       
                            (tmr_registers(0)(442) and tmr_registers(2)(442));                                                         
                                                                                                                                     
        global_tmr_voter(2)(443)  <=    (tmr_registers(0)(443) and tmr_registers(1)(443)) or                                            
                            (tmr_registers(1)(443) and tmr_registers(2)(443)) or                                                       
                            (tmr_registers(0)(443) and tmr_registers(2)(443));                                                         
                                                                                                                                     
        global_tmr_voter(2)(444)  <=    (tmr_registers(0)(444) and tmr_registers(1)(444)) or                                            
                            (tmr_registers(1)(444) and tmr_registers(2)(444)) or                                                       
                            (tmr_registers(0)(444) and tmr_registers(2)(444));                                                         
                                                                                                                                     
        global_tmr_voter(2)(445)  <=    (tmr_registers(0)(445) and tmr_registers(1)(445)) or                                            
                            (tmr_registers(1)(445) and tmr_registers(2)(445)) or                                                       
                            (tmr_registers(0)(445) and tmr_registers(2)(445));                                                         
                                                                                                                                     
        global_tmr_voter(2)(446)  <=    (tmr_registers(0)(446) and tmr_registers(1)(446)) or                                            
                            (tmr_registers(1)(446) and tmr_registers(2)(446)) or                                                       
                            (tmr_registers(0)(446) and tmr_registers(2)(446));                                                         
                                                                                                                                     
        global_tmr_voter(2)(447)  <=    (tmr_registers(0)(447) and tmr_registers(1)(447)) or                                            
                            (tmr_registers(1)(447) and tmr_registers(2)(447)) or                                                       
                            (tmr_registers(0)(447) and tmr_registers(2)(447));                                                         
                                                                                                                                     
        global_tmr_voter(2)(448)  <=    (tmr_registers(0)(448) and tmr_registers(1)(448)) or                                            
                            (tmr_registers(1)(448) and tmr_registers(2)(448)) or                                                       
                            (tmr_registers(0)(448) and tmr_registers(2)(448));                                                         
                                                                                                                                     
        global_tmr_voter(2)(449)  <=    (tmr_registers(0)(449) and tmr_registers(1)(449)) or                                            
                            (tmr_registers(1)(449) and tmr_registers(2)(449)) or                                                       
                            (tmr_registers(0)(449) and tmr_registers(2)(449));                                                         
                                                                                                                                     
        global_tmr_voter(2)(450)  <=    (tmr_registers(0)(450) and tmr_registers(1)(450)) or                                            
                            (tmr_registers(1)(450) and tmr_registers(2)(450)) or                                                       
                            (tmr_registers(0)(450) and tmr_registers(2)(450));                                                         
                                                                                                                                     
        global_tmr_voter(2)(451)  <=    (tmr_registers(0)(451) and tmr_registers(1)(451)) or                                            
                            (tmr_registers(1)(451) and tmr_registers(2)(451)) or                                                       
                            (tmr_registers(0)(451) and tmr_registers(2)(451));                                                         
                                                                                                                                     
        global_tmr_voter(2)(452)  <=    (tmr_registers(0)(452) and tmr_registers(1)(452)) or                                            
                            (tmr_registers(1)(452) and tmr_registers(2)(452)) or                                                       
                            (tmr_registers(0)(452) and tmr_registers(2)(452));                                                         
                                                                                                                                     
        global_tmr_voter(2)(453)  <=    (tmr_registers(0)(453) and tmr_registers(1)(453)) or                                            
                            (tmr_registers(1)(453) and tmr_registers(2)(453)) or                                                       
                            (tmr_registers(0)(453) and tmr_registers(2)(453));                                                         
                                                                                                                                     
        global_tmr_voter(2)(454)  <=    (tmr_registers(0)(454) and tmr_registers(1)(454)) or                                            
                            (tmr_registers(1)(454) and tmr_registers(2)(454)) or                                                       
                            (tmr_registers(0)(454) and tmr_registers(2)(454));                                                         
                                                                                                                                     
        global_tmr_voter(2)(455)  <=    (tmr_registers(0)(455) and tmr_registers(1)(455)) or                                            
                            (tmr_registers(1)(455) and tmr_registers(2)(455)) or                                                       
                            (tmr_registers(0)(455) and tmr_registers(2)(455));                                                         
                                                                                                                                     
        global_tmr_voter(2)(456)  <=    (tmr_registers(0)(456) and tmr_registers(1)(456)) or                                            
                            (tmr_registers(1)(456) and tmr_registers(2)(456)) or                                                       
                            (tmr_registers(0)(456) and tmr_registers(2)(456));                                                         
                                                                                                                                     
        global_tmr_voter(2)(457)  <=    (tmr_registers(0)(457) and tmr_registers(1)(457)) or                                            
                            (tmr_registers(1)(457) and tmr_registers(2)(457)) or                                                       
                            (tmr_registers(0)(457) and tmr_registers(2)(457));                                                         
                                                                                                                                     
        global_tmr_voter(2)(458)  <=    (tmr_registers(0)(458) and tmr_registers(1)(458)) or                                            
                            (tmr_registers(1)(458) and tmr_registers(2)(458)) or                                                       
                            (tmr_registers(0)(458) and tmr_registers(2)(458));                                                         
                                                                                                                                     
        global_tmr_voter(2)(459)  <=    (tmr_registers(0)(459) and tmr_registers(1)(459)) or                                            
                            (tmr_registers(1)(459) and tmr_registers(2)(459)) or                                                       
                            (tmr_registers(0)(459) and tmr_registers(2)(459));                                                         
                                                                                                                                     
        global_tmr_voter(2)(460)  <=    (tmr_registers(0)(460) and tmr_registers(1)(460)) or                                            
                            (tmr_registers(1)(460) and tmr_registers(2)(460)) or                                                       
                            (tmr_registers(0)(460) and tmr_registers(2)(460));                                                         
                                                                                                                                     
        global_tmr_voter(2)(461)  <=    (tmr_registers(0)(461) and tmr_registers(1)(461)) or                                            
                            (tmr_registers(1)(461) and tmr_registers(2)(461)) or                                                       
                            (tmr_registers(0)(461) and tmr_registers(2)(461));                                                         
                                                                                                                                     
        global_tmr_voter(2)(462)  <=    (tmr_registers(0)(462) and tmr_registers(1)(462)) or                                            
                            (tmr_registers(1)(462) and tmr_registers(2)(462)) or                                                       
                            (tmr_registers(0)(462) and tmr_registers(2)(462));                                                         
                                                                                                                                     
        global_tmr_voter(2)(463)  <=    (tmr_registers(0)(463) and tmr_registers(1)(463)) or                                            
                            (tmr_registers(1)(463) and tmr_registers(2)(463)) or                                                       
                            (tmr_registers(0)(463) and tmr_registers(2)(463));                                                         
                                                                                                                                     
        global_tmr_voter(2)(464)  <=    (tmr_registers(0)(464) and tmr_registers(1)(464)) or                                            
                            (tmr_registers(1)(464) and tmr_registers(2)(464)) or                                                       
                            (tmr_registers(0)(464) and tmr_registers(2)(464));                                                         
                                                                                                                                     
        global_tmr_voter(2)(465)  <=    (tmr_registers(0)(465) and tmr_registers(1)(465)) or                                            
                            (tmr_registers(1)(465) and tmr_registers(2)(465)) or                                                       
                            (tmr_registers(0)(465) and tmr_registers(2)(465));                                                         
                                                                                                                                     
        global_tmr_voter(2)(466)  <=    (tmr_registers(0)(466) and tmr_registers(1)(466)) or                                            
                            (tmr_registers(1)(466) and tmr_registers(2)(466)) or                                                       
                            (tmr_registers(0)(466) and tmr_registers(2)(466));                                                         
                                                                                                                                     
        global_tmr_voter(2)(467)  <=    (tmr_registers(0)(467) and tmr_registers(1)(467)) or                                            
                            (tmr_registers(1)(467) and tmr_registers(2)(467)) or                                                       
                            (tmr_registers(0)(467) and tmr_registers(2)(467));                                                         
                                                                                                                                     
        global_tmr_voter(2)(468)  <=    (tmr_registers(0)(468) and tmr_registers(1)(468)) or                                            
                            (tmr_registers(1)(468) and tmr_registers(2)(468)) or                                                       
                            (tmr_registers(0)(468) and tmr_registers(2)(468));                                                         
                                                                                                                                     
        global_tmr_voter(2)(469)  <=    (tmr_registers(0)(469) and tmr_registers(1)(469)) or                                            
                            (tmr_registers(1)(469) and tmr_registers(2)(469)) or                                                       
                            (tmr_registers(0)(469) and tmr_registers(2)(469));                                                         
                                                                                                                                     
        global_tmr_voter(2)(470)  <=    (tmr_registers(0)(470) and tmr_registers(1)(470)) or                                            
                            (tmr_registers(1)(470) and tmr_registers(2)(470)) or                                                       
                            (tmr_registers(0)(470) and tmr_registers(2)(470));                                                         
                                                                                                                                     
        global_tmr_voter(2)(471)  <=    (tmr_registers(0)(471) and tmr_registers(1)(471)) or                                            
                            (tmr_registers(1)(471) and tmr_registers(2)(471)) or                                                       
                            (tmr_registers(0)(471) and tmr_registers(2)(471));                                                         
                                                                                                                                     
        global_tmr_voter(2)(472)  <=    (tmr_registers(0)(472) and tmr_registers(1)(472)) or                                            
                            (tmr_registers(1)(472) and tmr_registers(2)(472)) or                                                       
                            (tmr_registers(0)(472) and tmr_registers(2)(472));                                                         
                                                                                                                                     
        global_tmr_voter(2)(473)  <=    (tmr_registers(0)(473) and tmr_registers(1)(473)) or                                            
                            (tmr_registers(1)(473) and tmr_registers(2)(473)) or                                                       
                            (tmr_registers(0)(473) and tmr_registers(2)(473));                                                         
                                                                                                                                     
        global_tmr_voter(2)(474)  <=    (tmr_registers(0)(474) and tmr_registers(1)(474)) or                                            
                            (tmr_registers(1)(474) and tmr_registers(2)(474)) or                                                       
                            (tmr_registers(0)(474) and tmr_registers(2)(474));                                                         
                                                                                                                                     
        global_tmr_voter(2)(475)  <=    (tmr_registers(0)(475) and tmr_registers(1)(475)) or                                            
                            (tmr_registers(1)(475) and tmr_registers(2)(475)) or                                                       
                            (tmr_registers(0)(475) and tmr_registers(2)(475));                                                         
                                                                                                                                     
        global_tmr_voter(2)(476)  <=    (tmr_registers(0)(476) and tmr_registers(1)(476)) or                                            
                            (tmr_registers(1)(476) and tmr_registers(2)(476)) or                                                       
                            (tmr_registers(0)(476) and tmr_registers(2)(476));                                                         
                                                                                                                                     
        global_tmr_voter(2)(477)  <=    (tmr_registers(0)(477) and tmr_registers(1)(477)) or                                            
                            (tmr_registers(1)(477) and tmr_registers(2)(477)) or                                                       
                            (tmr_registers(0)(477) and tmr_registers(2)(477));                                                         
                                                                                                                                     
        global_tmr_voter(2)(478)  <=    (tmr_registers(0)(478) and tmr_registers(1)(478)) or                                            
                            (tmr_registers(1)(478) and tmr_registers(2)(478)) or                                                       
                            (tmr_registers(0)(478) and tmr_registers(2)(478));                                                         
                                                                                                                                     
        global_tmr_voter(2)(479)  <=    (tmr_registers(0)(479) and tmr_registers(1)(479)) or                                            
                            (tmr_registers(1)(479) and tmr_registers(2)(479)) or                                                       
                            (tmr_registers(0)(479) and tmr_registers(2)(479));                                                         
                                                                                                                                     
        global_tmr_voter(2)(480)  <=    (tmr_registers(0)(480) and tmr_registers(1)(480)) or                                            
                            (tmr_registers(1)(480) and tmr_registers(2)(480)) or                                                       
                            (tmr_registers(0)(480) and tmr_registers(2)(480));                                                         
                                                                                                                                     
        global_tmr_voter(2)(481)  <=    (tmr_registers(0)(481) and tmr_registers(1)(481)) or                                            
                            (tmr_registers(1)(481) and tmr_registers(2)(481)) or                                                       
                            (tmr_registers(0)(481) and tmr_registers(2)(481));                                                         
                                                                                                                                     
        global_tmr_voter(2)(482)  <=    (tmr_registers(0)(482) and tmr_registers(1)(482)) or                                            
                            (tmr_registers(1)(482) and tmr_registers(2)(482)) or                                                       
                            (tmr_registers(0)(482) and tmr_registers(2)(482));                                                         
                                                                                                                                     
        global_tmr_voter(2)(483)  <=    (tmr_registers(0)(483) and tmr_registers(1)(483)) or                                            
                            (tmr_registers(1)(483) and tmr_registers(2)(483)) or                                                       
                            (tmr_registers(0)(483) and tmr_registers(2)(483));                                                         
                                                                                                                                     
        global_tmr_voter(2)(484)  <=    (tmr_registers(0)(484) and tmr_registers(1)(484)) or                                            
                            (tmr_registers(1)(484) and tmr_registers(2)(484)) or                                                       
                            (tmr_registers(0)(484) and tmr_registers(2)(484));                                                         
                                                                                                                                     
        global_tmr_voter(2)(485)  <=    (tmr_registers(0)(485) and tmr_registers(1)(485)) or                                            
                            (tmr_registers(1)(485) and tmr_registers(2)(485)) or                                                       
                            (tmr_registers(0)(485) and tmr_registers(2)(485));                                                         
                                                                                                                                     
        global_tmr_voter(2)(486)  <=    (tmr_registers(0)(486) and tmr_registers(1)(486)) or                                            
                            (tmr_registers(1)(486) and tmr_registers(2)(486)) or                                                       
                            (tmr_registers(0)(486) and tmr_registers(2)(486));                                                         
                                                                                                                                     
        global_tmr_voter(2)(487)  <=    (tmr_registers(0)(487) and tmr_registers(1)(487)) or                                            
                            (tmr_registers(1)(487) and tmr_registers(2)(487)) or                                                       
                            (tmr_registers(0)(487) and tmr_registers(2)(487));                                                         
                                                                                                                                     
        global_tmr_voter(2)(488)  <=    (tmr_registers(0)(488) and tmr_registers(1)(488)) or                                            
                            (tmr_registers(1)(488) and tmr_registers(2)(488)) or                                                       
                            (tmr_registers(0)(488) and tmr_registers(2)(488));                                                         
                                                                                                                                     
        global_tmr_voter(2)(489)  <=    (tmr_registers(0)(489) and tmr_registers(1)(489)) or                                            
                            (tmr_registers(1)(489) and tmr_registers(2)(489)) or                                                       
                            (tmr_registers(0)(489) and tmr_registers(2)(489));                                                         
                                                                                                                                     
        global_tmr_voter(2)(490)  <=    (tmr_registers(0)(490) and tmr_registers(1)(490)) or                                            
                            (tmr_registers(1)(490) and tmr_registers(2)(490)) or                                                       
                            (tmr_registers(0)(490) and tmr_registers(2)(490));                                                         
                                                                                                                                     
        global_tmr_voter(2)(491)  <=    (tmr_registers(0)(491) and tmr_registers(1)(491)) or                                            
                            (tmr_registers(1)(491) and tmr_registers(2)(491)) or                                                       
                            (tmr_registers(0)(491) and tmr_registers(2)(491));                                                         
                                                                                                                                     
        global_tmr_voter(2)(492)  <=    (tmr_registers(0)(492) and tmr_registers(1)(492)) or                                            
                            (tmr_registers(1)(492) and tmr_registers(2)(492)) or                                                       
                            (tmr_registers(0)(492) and tmr_registers(2)(492));                                                         
                                                                                                                                     
        global_tmr_voter(2)(493)  <=    (tmr_registers(0)(493) and tmr_registers(1)(493)) or                                            
                            (tmr_registers(1)(493) and tmr_registers(2)(493)) or                                                       
                            (tmr_registers(0)(493) and tmr_registers(2)(493));                                                         
                                                                                                                                     
        global_tmr_voter(2)(494)  <=    (tmr_registers(0)(494) and tmr_registers(1)(494)) or                                            
                            (tmr_registers(1)(494) and tmr_registers(2)(494)) or                                                       
                            (tmr_registers(0)(494) and tmr_registers(2)(494));                                                         
                                                                                                                                     
        global_tmr_voter(2)(495)  <=    (tmr_registers(0)(495) and tmr_registers(1)(495)) or                                            
                            (tmr_registers(1)(495) and tmr_registers(2)(495)) or                                                       
                            (tmr_registers(0)(495) and tmr_registers(2)(495));                                                         
                                                                                                                                     
        global_tmr_voter(2)(496)  <=    (tmr_registers(0)(496) and tmr_registers(1)(496)) or                                            
                            (tmr_registers(1)(496) and tmr_registers(2)(496)) or                                                       
                            (tmr_registers(0)(496) and tmr_registers(2)(496));                                                         
                                                                                                                                     
        global_tmr_voter(2)(497)  <=    (tmr_registers(0)(497) and tmr_registers(1)(497)) or                                            
                            (tmr_registers(1)(497) and tmr_registers(2)(497)) or                                                       
                            (tmr_registers(0)(497) and tmr_registers(2)(497));                                                         
                                                                                                                                     
        global_tmr_voter(2)(498)  <=    (tmr_registers(0)(498) and tmr_registers(1)(498)) or                                            
                            (tmr_registers(1)(498) and tmr_registers(2)(498)) or                                                       
                            (tmr_registers(0)(498) and tmr_registers(2)(498));                                                         
                                                                                                                                     
        global_tmr_voter(2)(499)  <=    (tmr_registers(0)(499) and tmr_registers(1)(499)) or                                            
                            (tmr_registers(1)(499) and tmr_registers(2)(499)) or                                                       
                            (tmr_registers(0)(499) and tmr_registers(2)(499));                                                         
                                                                                                                                     
        global_tmr_voter(2)(500)  <=    (tmr_registers(0)(500) and tmr_registers(1)(500)) or                                            
                            (tmr_registers(1)(500) and tmr_registers(2)(500)) or                                                       
                            (tmr_registers(0)(500) and tmr_registers(2)(500));                                                         
                                                                                                                                     
        global_tmr_voter(2)(501)  <=    (tmr_registers(0)(501) and tmr_registers(1)(501)) or                                            
                            (tmr_registers(1)(501) and tmr_registers(2)(501)) or                                                       
                            (tmr_registers(0)(501) and tmr_registers(2)(501));                                                         
                                                                                                                                     
        global_tmr_voter(2)(502)  <=    (tmr_registers(0)(502) and tmr_registers(1)(502)) or                                            
                            (tmr_registers(1)(502) and tmr_registers(2)(502)) or                                                       
                            (tmr_registers(0)(502) and tmr_registers(2)(502));                                                         
                                                                                                                                     
        global_tmr_voter(2)(503)  <=    (tmr_registers(0)(503) and tmr_registers(1)(503)) or                                            
                            (tmr_registers(1)(503) and tmr_registers(2)(503)) or                                                       
                            (tmr_registers(0)(503) and tmr_registers(2)(503));                                                         
                                                                                                                                     
        global_tmr_voter(2)(504)  <=    (tmr_registers(0)(504) and tmr_registers(1)(504)) or                                            
                            (tmr_registers(1)(504) and tmr_registers(2)(504)) or                                                       
                            (tmr_registers(0)(504) and tmr_registers(2)(504));                                                         
                                                                                                                                     
        global_tmr_voter(2)(505)  <=    (tmr_registers(0)(505) and tmr_registers(1)(505)) or                                            
                            (tmr_registers(1)(505) and tmr_registers(2)(505)) or                                                       
                            (tmr_registers(0)(505) and tmr_registers(2)(505));                                                         
                                                                                                                                     
        global_tmr_voter(2)(506)  <=    (tmr_registers(0)(506) and tmr_registers(1)(506)) or                                            
                            (tmr_registers(1)(506) and tmr_registers(2)(506)) or                                                       
                            (tmr_registers(0)(506) and tmr_registers(2)(506));                                                         
                                                                                                                                     
        global_tmr_voter(2)(507)  <=    (tmr_registers(0)(507) and tmr_registers(1)(507)) or                                            
                            (tmr_registers(1)(507) and tmr_registers(2)(507)) or                                                       
                            (tmr_registers(0)(507) and tmr_registers(2)(507));                                                         
                                                                                                                                     
        global_tmr_voter(2)(508)  <=    (tmr_registers(0)(508) and tmr_registers(1)(508)) or                                            
                            (tmr_registers(1)(508) and tmr_registers(2)(508)) or                                                       
                            (tmr_registers(0)(508) and tmr_registers(2)(508));                                                         
                                                                                                                                     
        global_tmr_voter(2)(509)  <=    (tmr_registers(0)(509) and tmr_registers(1)(509)) or                                            
                            (tmr_registers(1)(509) and tmr_registers(2)(509)) or                                                       
                            (tmr_registers(0)(509) and tmr_registers(2)(509));                                                         
                                                                                                                                     
        global_tmr_voter(2)(510)  <=    (tmr_registers(0)(510) and tmr_registers(1)(510)) or                                            
                            (tmr_registers(1)(510) and tmr_registers(2)(510)) or                                                       
                            (tmr_registers(0)(510) and tmr_registers(2)(510));                                                         
                                                                                                                                     
        global_tmr_voter(2)(511)  <=    (tmr_registers(0)(511) and tmr_registers(1)(511)) or                                            
                            (tmr_registers(1)(511) and tmr_registers(2)(511)) or                                                       
                            (tmr_registers(0)(511) and tmr_registers(2)(511));                                                         
                                                                                                                                     
        global_tmr_voter(2)(512)  <=    (tmr_registers(0)(512) and tmr_registers(1)(512)) or                                            
                            (tmr_registers(1)(512) and tmr_registers(2)(512)) or                                                       
                            (tmr_registers(0)(512) and tmr_registers(2)(512));                                                         
                                                                                                                                     
        global_tmr_voter(2)(513)  <=    (tmr_registers(0)(513) and tmr_registers(1)(513)) or                                            
                            (tmr_registers(1)(513) and tmr_registers(2)(513)) or                                                       
                            (tmr_registers(0)(513) and tmr_registers(2)(513));                                                         
                                                                                                                                     
        global_tmr_voter(2)(514)  <=    (tmr_registers(0)(514) and tmr_registers(1)(514)) or                                            
                            (tmr_registers(1)(514) and tmr_registers(2)(514)) or                                                       
                            (tmr_registers(0)(514) and tmr_registers(2)(514));                                                         
                                                                                                                                     
        global_tmr_voter(2)(515)  <=    (tmr_registers(0)(515) and tmr_registers(1)(515)) or                                            
                            (tmr_registers(1)(515) and tmr_registers(2)(515)) or                                                       
                            (tmr_registers(0)(515) and tmr_registers(2)(515));                                                         
                                                                                                                                     
        global_tmr_voter(2)(516)  <=    (tmr_registers(0)(516) and tmr_registers(1)(516)) or                                            
                            (tmr_registers(1)(516) and tmr_registers(2)(516)) or                                                       
                            (tmr_registers(0)(516) and tmr_registers(2)(516));                                                         
                                                                                                                                     
        global_tmr_voter(2)(517)  <=    (tmr_registers(0)(517) and tmr_registers(1)(517)) or                                            
                            (tmr_registers(1)(517) and tmr_registers(2)(517)) or                                                       
                            (tmr_registers(0)(517) and tmr_registers(2)(517));                                                         
                                                                                                                                     
        global_tmr_voter(2)(518)  <=    (tmr_registers(0)(518) and tmr_registers(1)(518)) or                                            
                            (tmr_registers(1)(518) and tmr_registers(2)(518)) or                                                       
                            (tmr_registers(0)(518) and tmr_registers(2)(518));                                                         
                                                                                                                                     
        global_tmr_voter(2)(519)  <=    (tmr_registers(0)(519) and tmr_registers(1)(519)) or                                            
                            (tmr_registers(1)(519) and tmr_registers(2)(519)) or                                                       
                            (tmr_registers(0)(519) and tmr_registers(2)(519));                                                         
                                                                                                                                     
        global_tmr_voter(2)(520)  <=    (tmr_registers(0)(520) and tmr_registers(1)(520)) or                                            
                            (tmr_registers(1)(520) and tmr_registers(2)(520)) or                                                       
                            (tmr_registers(0)(520) and tmr_registers(2)(520));                                                         
                                                                                                                                     
        global_tmr_voter(2)(521)  <=    (tmr_registers(0)(521) and tmr_registers(1)(521)) or                                            
                            (tmr_registers(1)(521) and tmr_registers(2)(521)) or                                                       
                            (tmr_registers(0)(521) and tmr_registers(2)(521));                                                         
                                                                                                                                     
        global_tmr_voter(2)(522)  <=    (tmr_registers(0)(522) and tmr_registers(1)(522)) or                                            
                            (tmr_registers(1)(522) and tmr_registers(2)(522)) or                                                       
                            (tmr_registers(0)(522) and tmr_registers(2)(522));                                                         
                                                                                                                                     
        global_tmr_voter(2)(523)  <=    (tmr_registers(0)(523) and tmr_registers(1)(523)) or                                            
                            (tmr_registers(1)(523) and tmr_registers(2)(523)) or                                                       
                            (tmr_registers(0)(523) and tmr_registers(2)(523));                                                         
                                                                                                                                     
        global_tmr_voter(2)(524)  <=    (tmr_registers(0)(524) and tmr_registers(1)(524)) or                                            
                            (tmr_registers(1)(524) and tmr_registers(2)(524)) or                                                       
                            (tmr_registers(0)(524) and tmr_registers(2)(524));                                                         
                                                                                                                                     
        global_tmr_voter(2)(525)  <=    (tmr_registers(0)(525) and tmr_registers(1)(525)) or                                            
                            (tmr_registers(1)(525) and tmr_registers(2)(525)) or                                                       
                            (tmr_registers(0)(525) and tmr_registers(2)(525));                                                         
                                                                                                                                     
        global_tmr_voter(2)(526)  <=    (tmr_registers(0)(526) and tmr_registers(1)(526)) or                                            
                            (tmr_registers(1)(526) and tmr_registers(2)(526)) or                                                       
                            (tmr_registers(0)(526) and tmr_registers(2)(526));                                                         
                                                                                                                                     
        global_tmr_voter(2)(527)  <=    (tmr_registers(0)(527) and tmr_registers(1)(527)) or                                            
                            (tmr_registers(1)(527) and tmr_registers(2)(527)) or                                                       
                            (tmr_registers(0)(527) and tmr_registers(2)(527));                                                         
                                                                                                                                     
        global_tmr_voter(2)(528)  <=    (tmr_registers(0)(528) and tmr_registers(1)(528)) or                                            
                            (tmr_registers(1)(528) and tmr_registers(2)(528)) or                                                       
                            (tmr_registers(0)(528) and tmr_registers(2)(528));                                                         
                                                                                                                                     
        global_tmr_voter(2)(529)  <=    (tmr_registers(0)(529) and tmr_registers(1)(529)) or                                            
                            (tmr_registers(1)(529) and tmr_registers(2)(529)) or                                                       
                            (tmr_registers(0)(529) and tmr_registers(2)(529));                                                         
                                                                                                                                     
        global_tmr_voter(2)(530)  <=    (tmr_registers(0)(530) and tmr_registers(1)(530)) or                                            
                            (tmr_registers(1)(530) and tmr_registers(2)(530)) or                                                       
                            (tmr_registers(0)(530) and tmr_registers(2)(530));                                                         
                                                                                                                                     
        global_tmr_voter(2)(531)  <=    (tmr_registers(0)(531) and tmr_registers(1)(531)) or                                            
                            (tmr_registers(1)(531) and tmr_registers(2)(531)) or                                                       
                            (tmr_registers(0)(531) and tmr_registers(2)(531));                                                         
                                                                                                                                     
        global_tmr_voter(2)(532)  <=    (tmr_registers(0)(532) and tmr_registers(1)(532)) or                                            
                            (tmr_registers(1)(532) and tmr_registers(2)(532)) or                                                       
                            (tmr_registers(0)(532) and tmr_registers(2)(532));                                                         
                                                                                                                                     
        global_tmr_voter(2)(533)  <=    (tmr_registers(0)(533) and tmr_registers(1)(533)) or                                            
                            (tmr_registers(1)(533) and tmr_registers(2)(533)) or                                                       
                            (tmr_registers(0)(533) and tmr_registers(2)(533));                                                         
                                                                                                                                     
        global_tmr_voter(2)(534)  <=    (tmr_registers(0)(534) and tmr_registers(1)(534)) or                                            
                            (tmr_registers(1)(534) and tmr_registers(2)(534)) or                                                       
                            (tmr_registers(0)(534) and tmr_registers(2)(534));                                                         
                                                                                                                                     
        global_tmr_voter(2)(535)  <=    (tmr_registers(0)(535) and tmr_registers(1)(535)) or                                            
                            (tmr_registers(1)(535) and tmr_registers(2)(535)) or                                                       
                            (tmr_registers(0)(535) and tmr_registers(2)(535));                                                         
                                                                                                                                     
        global_tmr_voter(2)(536)  <=    (tmr_registers(0)(536) and tmr_registers(1)(536)) or                                            
                            (tmr_registers(1)(536) and tmr_registers(2)(536)) or                                                       
                            (tmr_registers(0)(536) and tmr_registers(2)(536));                                                         
                                                                                                                                     
        global_tmr_voter(2)(537)  <=    (tmr_registers(0)(537) and tmr_registers(1)(537)) or                                            
                            (tmr_registers(1)(537) and tmr_registers(2)(537)) or                                                       
                            (tmr_registers(0)(537) and tmr_registers(2)(537));                                                         
                                                                                                                                     
        global_tmr_voter(2)(538)  <=    (tmr_registers(0)(538) and tmr_registers(1)(538)) or                                            
                            (tmr_registers(1)(538) and tmr_registers(2)(538)) or                                                       
                            (tmr_registers(0)(538) and tmr_registers(2)(538));                                                         
                                                                                                                                     
        global_tmr_voter(2)(539)  <=    (tmr_registers(0)(539) and tmr_registers(1)(539)) or                                            
                            (tmr_registers(1)(539) and tmr_registers(2)(539)) or                                                       
                            (tmr_registers(0)(539) and tmr_registers(2)(539));                                                         
                                                                                                                                     
        global_tmr_voter(2)(540)  <=    (tmr_registers(0)(540) and tmr_registers(1)(540)) or                                            
                            (tmr_registers(1)(540) and tmr_registers(2)(540)) or                                                       
                            (tmr_registers(0)(540) and tmr_registers(2)(540));                                                         
                                                                                                                                     
        global_tmr_voter(2)(541)  <=    (tmr_registers(0)(541) and tmr_registers(1)(541)) or                                            
                            (tmr_registers(1)(541) and tmr_registers(2)(541)) or                                                       
                            (tmr_registers(0)(541) and tmr_registers(2)(541));                                                         
                                                                                                                                     
        global_tmr_voter(2)(542)  <=    (tmr_registers(0)(542) and tmr_registers(1)(542)) or                                            
                            (tmr_registers(1)(542) and tmr_registers(2)(542)) or                                                       
                            (tmr_registers(0)(542) and tmr_registers(2)(542));                                                         
                                                                                                                                     
        global_tmr_voter(2)(543)  <=    (tmr_registers(0)(543) and tmr_registers(1)(543)) or                                            
                            (tmr_registers(1)(543) and tmr_registers(2)(543)) or                                                       
                            (tmr_registers(0)(543) and tmr_registers(2)(543));                                                         
                                                                                                                                     
        global_tmr_voter(2)(544)  <=    (tmr_registers(0)(544) and tmr_registers(1)(544)) or                                            
                            (tmr_registers(1)(544) and tmr_registers(2)(544)) or                                                       
                            (tmr_registers(0)(544) and tmr_registers(2)(544));                                                         
                                                                                                                                     
        global_tmr_voter(2)(545)  <=    (tmr_registers(0)(545) and tmr_registers(1)(545)) or                                            
                            (tmr_registers(1)(545) and tmr_registers(2)(545)) or                                                       
                            (tmr_registers(0)(545) and tmr_registers(2)(545));                                                         
                                                                                                                                     
        global_tmr_voter(2)(546)  <=    (tmr_registers(0)(546) and tmr_registers(1)(546)) or                                            
                            (tmr_registers(1)(546) and tmr_registers(2)(546)) or                                                       
                            (tmr_registers(0)(546) and tmr_registers(2)(546));                                                         
                                                                                                                                     
        global_tmr_voter(2)(547)  <=    (tmr_registers(0)(547) and tmr_registers(1)(547)) or                                            
                            (tmr_registers(1)(547) and tmr_registers(2)(547)) or                                                       
                            (tmr_registers(0)(547) and tmr_registers(2)(547));                                                         
                                                                                                                                     
        global_tmr_voter(2)(548)  <=    (tmr_registers(0)(548) and tmr_registers(1)(548)) or                                            
                            (tmr_registers(1)(548) and tmr_registers(2)(548)) or                                                       
                            (tmr_registers(0)(548) and tmr_registers(2)(548));                                                         
                                                                                                                                     
        global_tmr_voter(2)(549)  <=    (tmr_registers(0)(549) and tmr_registers(1)(549)) or                                            
                            (tmr_registers(1)(549) and tmr_registers(2)(549)) or                                                       
                            (tmr_registers(0)(549) and tmr_registers(2)(549));                                                         
                                                                                                                                     
        global_tmr_voter(2)(550)  <=    (tmr_registers(0)(550) and tmr_registers(1)(550)) or                                            
                            (tmr_registers(1)(550) and tmr_registers(2)(550)) or                                                       
                            (tmr_registers(0)(550) and tmr_registers(2)(550));                                                         
                                                                                                                                     
        global_tmr_voter(2)(551)  <=    (tmr_registers(0)(551) and tmr_registers(1)(551)) or                                            
                            (tmr_registers(1)(551) and tmr_registers(2)(551)) or                                                       
                            (tmr_registers(0)(551) and tmr_registers(2)(551));                                                         
                                                                                                                                     
        global_tmr_voter(2)(552)  <=    (tmr_registers(0)(552) and tmr_registers(1)(552)) or                                            
                            (tmr_registers(1)(552) and tmr_registers(2)(552)) or                                                       
                            (tmr_registers(0)(552) and tmr_registers(2)(552));                                                         
                                                                                                                                     
        global_tmr_voter(2)(553)  <=    (tmr_registers(0)(553) and tmr_registers(1)(553)) or                                            
                            (tmr_registers(1)(553) and tmr_registers(2)(553)) or                                                       
                            (tmr_registers(0)(553) and tmr_registers(2)(553));                                                         
                                                                                                                                     
        global_tmr_voter(2)(554)  <=    (tmr_registers(0)(554) and tmr_registers(1)(554)) or                                            
                            (tmr_registers(1)(554) and tmr_registers(2)(554)) or                                                       
                            (tmr_registers(0)(554) and tmr_registers(2)(554));                                                         
                                                                                                                                     
        global_tmr_voter(2)(555)  <=    (tmr_registers(0)(555) and tmr_registers(1)(555)) or                                            
                            (tmr_registers(1)(555) and tmr_registers(2)(555)) or                                                       
                            (tmr_registers(0)(555) and tmr_registers(2)(555));                                                         
                                                                                                                                     
        global_tmr_voter(2)(556)  <=    (tmr_registers(0)(556) and tmr_registers(1)(556)) or                                            
                            (tmr_registers(1)(556) and tmr_registers(2)(556)) or                                                       
                            (tmr_registers(0)(556) and tmr_registers(2)(556));                                                         
                                                                                                                                     
        global_tmr_voter(2)(557)  <=    (tmr_registers(0)(557) and tmr_registers(1)(557)) or                                            
                            (tmr_registers(1)(557) and tmr_registers(2)(557)) or                                                       
                            (tmr_registers(0)(557) and tmr_registers(2)(557));                                                         
                                                                                                                                     
        global_tmr_voter(2)(558)  <=    (tmr_registers(0)(558) and tmr_registers(1)(558)) or                                            
                            (tmr_registers(1)(558) and tmr_registers(2)(558)) or                                                       
                            (tmr_registers(0)(558) and tmr_registers(2)(558));                                                         
                                                                                                                                     
        global_tmr_voter(2)(559)  <=    (tmr_registers(0)(559) and tmr_registers(1)(559)) or                                            
                            (tmr_registers(1)(559) and tmr_registers(2)(559)) or                                                       
                            (tmr_registers(0)(559) and tmr_registers(2)(559));                                                         
                                                                                                                                     
        global_tmr_voter(2)(560)  <=    (tmr_registers(0)(560) and tmr_registers(1)(560)) or                                            
                            (tmr_registers(1)(560) and tmr_registers(2)(560)) or                                                       
                            (tmr_registers(0)(560) and tmr_registers(2)(560));                                                         
                                                                                                                                     
        global_tmr_voter(2)(561)  <=    (tmr_registers(0)(561) and tmr_registers(1)(561)) or                                            
                            (tmr_registers(1)(561) and tmr_registers(2)(561)) or                                                       
                            (tmr_registers(0)(561) and tmr_registers(2)(561));                                                         
                                                                                                                                     
        global_tmr_voter(2)(562)  <=    (tmr_registers(0)(562) and tmr_registers(1)(562)) or                                            
                            (tmr_registers(1)(562) and tmr_registers(2)(562)) or                                                       
                            (tmr_registers(0)(562) and tmr_registers(2)(562));                                                         
                                                                                                                                     
        global_tmr_voter(2)(563)  <=    (tmr_registers(0)(563) and tmr_registers(1)(563)) or                                            
                            (tmr_registers(1)(563) and tmr_registers(2)(563)) or                                                       
                            (tmr_registers(0)(563) and tmr_registers(2)(563));                                                         
                                                                                                                                     
        global_tmr_voter(2)(564)  <=    (tmr_registers(0)(564) and tmr_registers(1)(564)) or                                            
                            (tmr_registers(1)(564) and tmr_registers(2)(564)) or                                                       
                            (tmr_registers(0)(564) and tmr_registers(2)(564));                                                         
                                                                                                                                     
        global_tmr_voter(2)(565)  <=    (tmr_registers(0)(565) and tmr_registers(1)(565)) or                                            
                            (tmr_registers(1)(565) and tmr_registers(2)(565)) or                                                       
                            (tmr_registers(0)(565) and tmr_registers(2)(565));                                                         
                                                                                                                                     
        global_tmr_voter(2)(566)  <=    (tmr_registers(0)(566) and tmr_registers(1)(566)) or                                            
                            (tmr_registers(1)(566) and tmr_registers(2)(566)) or                                                       
                            (tmr_registers(0)(566) and tmr_registers(2)(566));                                                         
                                                                                                                                     
        global_tmr_voter(2)(567)  <=    (tmr_registers(0)(567) and tmr_registers(1)(567)) or                                            
                            (tmr_registers(1)(567) and tmr_registers(2)(567)) or                                                       
                            (tmr_registers(0)(567) and tmr_registers(2)(567));                                                         
                                                                                                                                     
        global_tmr_voter(2)(568)  <=    (tmr_registers(0)(568) and tmr_registers(1)(568)) or                                            
                            (tmr_registers(1)(568) and tmr_registers(2)(568)) or                                                       
                            (tmr_registers(0)(568) and tmr_registers(2)(568));                                                         
                                                                                                                                     
        global_tmr_voter(2)(569)  <=    (tmr_registers(0)(569) and tmr_registers(1)(569)) or                                            
                            (tmr_registers(1)(569) and tmr_registers(2)(569)) or                                                       
                            (tmr_registers(0)(569) and tmr_registers(2)(569));                                                         
                                                                                                                                     
        global_tmr_voter(2)(570)  <=    (tmr_registers(0)(570) and tmr_registers(1)(570)) or                                            
                            (tmr_registers(1)(570) and tmr_registers(2)(570)) or                                                       
                            (tmr_registers(0)(570) and tmr_registers(2)(570));                                                         
                                                                                                                                     
        global_tmr_voter(2)(571)  <=    (tmr_registers(0)(571) and tmr_registers(1)(571)) or                                            
                            (tmr_registers(1)(571) and tmr_registers(2)(571)) or                                                       
                            (tmr_registers(0)(571) and tmr_registers(2)(571));                                                         
                                                                                                                                     
        global_tmr_voter(2)(572)  <=    (tmr_registers(0)(572) and tmr_registers(1)(572)) or                                            
                            (tmr_registers(1)(572) and tmr_registers(2)(572)) or                                                       
                            (tmr_registers(0)(572) and tmr_registers(2)(572));                                                         
                                                                                                                                     
        global_tmr_voter(2)(573)  <=    (tmr_registers(0)(573) and tmr_registers(1)(573)) or                                            
                            (tmr_registers(1)(573) and tmr_registers(2)(573)) or                                                       
                            (tmr_registers(0)(573) and tmr_registers(2)(573));                                                         
                                                                                                                                     
        global_tmr_voter(2)(574)  <=    (tmr_registers(0)(574) and tmr_registers(1)(574)) or                                            
                            (tmr_registers(1)(574) and tmr_registers(2)(574)) or                                                       
                            (tmr_registers(0)(574) and tmr_registers(2)(574));                                                         
                                                                                                                                     
        global_tmr_voter(2)(575)  <=    (tmr_registers(0)(575) and tmr_registers(1)(575)) or                                            
                            (tmr_registers(1)(575) and tmr_registers(2)(575)) or                                                       
                            (tmr_registers(0)(575) and tmr_registers(2)(575));                                                         
                                                                                                                                     
        global_tmr_voter(2)(576)  <=    (tmr_registers(0)(576) and tmr_registers(1)(576)) or                                            
                            (tmr_registers(1)(576) and tmr_registers(2)(576)) or                                                       
                            (tmr_registers(0)(576) and tmr_registers(2)(576));                                                         
                                                                                                                                     
        global_tmr_voter(2)(577)  <=    (tmr_registers(0)(577) and tmr_registers(1)(577)) or                                            
                            (tmr_registers(1)(577) and tmr_registers(2)(577)) or                                                       
                            (tmr_registers(0)(577) and tmr_registers(2)(577));                                                         
                                                                                                                                     
        global_tmr_voter(2)(578)  <=    (tmr_registers(0)(578) and tmr_registers(1)(578)) or                                            
                            (tmr_registers(1)(578) and tmr_registers(2)(578)) or                                                       
                            (tmr_registers(0)(578) and tmr_registers(2)(578));                                                         
                                                                                                                                     
        global_tmr_voter(2)(579)  <=    (tmr_registers(0)(579) and tmr_registers(1)(579)) or                                            
                            (tmr_registers(1)(579) and tmr_registers(2)(579)) or                                                       
                            (tmr_registers(0)(579) and tmr_registers(2)(579));                                                         
                                                                                                                                     
        global_tmr_voter(2)(580)  <=    (tmr_registers(0)(580) and tmr_registers(1)(580)) or                                            
                            (tmr_registers(1)(580) and tmr_registers(2)(580)) or                                                       
                            (tmr_registers(0)(580) and tmr_registers(2)(580));                                                         
                                                                                                                                     
        global_tmr_voter(2)(581)  <=    (tmr_registers(0)(581) and tmr_registers(1)(581)) or                                            
                            (tmr_registers(1)(581) and tmr_registers(2)(581)) or                                                       
                            (tmr_registers(0)(581) and tmr_registers(2)(581));                                                         
                                                                                                                                     
        global_tmr_voter(2)(582)  <=    (tmr_registers(0)(582) and tmr_registers(1)(582)) or                                            
                            (tmr_registers(1)(582) and tmr_registers(2)(582)) or                                                       
                            (tmr_registers(0)(582) and tmr_registers(2)(582));                                                         
                                                                                                                                     
        global_tmr_voter(2)(583)  <=    (tmr_registers(0)(583) and tmr_registers(1)(583)) or                                            
                            (tmr_registers(1)(583) and tmr_registers(2)(583)) or                                                       
                            (tmr_registers(0)(583) and tmr_registers(2)(583));                                                         
                                                                                                                                     
        global_tmr_voter(2)(584)  <=    (tmr_registers(0)(584) and tmr_registers(1)(584)) or                                            
                            (tmr_registers(1)(584) and tmr_registers(2)(584)) or                                                       
                            (tmr_registers(0)(584) and tmr_registers(2)(584));                                                         
                                                                                                                                     
        global_tmr_voter(2)(585)  <=    (tmr_registers(0)(585) and tmr_registers(1)(585)) or                                            
                            (tmr_registers(1)(585) and tmr_registers(2)(585)) or                                                       
                            (tmr_registers(0)(585) and tmr_registers(2)(585));                                                         
                                                                                                                                     
        global_tmr_voter(2)(586)  <=    (tmr_registers(0)(586) and tmr_registers(1)(586)) or                                            
                            (tmr_registers(1)(586) and tmr_registers(2)(586)) or                                                       
                            (tmr_registers(0)(586) and tmr_registers(2)(586));                                                         
                                                                                                                                     
        global_tmr_voter(2)(587)  <=    (tmr_registers(0)(587) and tmr_registers(1)(587)) or                                            
                            (tmr_registers(1)(587) and tmr_registers(2)(587)) or                                                       
                            (tmr_registers(0)(587) and tmr_registers(2)(587));                                                         
                                                                                                                                     
        global_tmr_voter(2)(588)  <=    (tmr_registers(0)(588) and tmr_registers(1)(588)) or                                            
                            (tmr_registers(1)(588) and tmr_registers(2)(588)) or                                                       
                            (tmr_registers(0)(588) and tmr_registers(2)(588));                                                         
                                                                                                                                     
        global_tmr_voter(2)(589)  <=    (tmr_registers(0)(589) and tmr_registers(1)(589)) or                                            
                            (tmr_registers(1)(589) and tmr_registers(2)(589)) or                                                       
                            (tmr_registers(0)(589) and tmr_registers(2)(589));                                                         
                                                                                                                                     
        global_tmr_voter(2)(590)  <=    (tmr_registers(0)(590) and tmr_registers(1)(590)) or                                            
                            (tmr_registers(1)(590) and tmr_registers(2)(590)) or                                                       
                            (tmr_registers(0)(590) and tmr_registers(2)(590));                                                         
                                                                                                                                     
        global_tmr_voter(2)(591)  <=    (tmr_registers(0)(591) and tmr_registers(1)(591)) or                                            
                            (tmr_registers(1)(591) and tmr_registers(2)(591)) or                                                       
                            (tmr_registers(0)(591) and tmr_registers(2)(591));                                                         
                                                                                                                                     
        global_tmr_voter(2)(592)  <=    (tmr_registers(0)(592) and tmr_registers(1)(592)) or                                            
                            (tmr_registers(1)(592) and tmr_registers(2)(592)) or                                                       
                            (tmr_registers(0)(592) and tmr_registers(2)(592));                                                         
                                                                                                                                     
        global_tmr_voter(2)(593)  <=    (tmr_registers(0)(593) and tmr_registers(1)(593)) or                                            
                            (tmr_registers(1)(593) and tmr_registers(2)(593)) or                                                       
                            (tmr_registers(0)(593) and tmr_registers(2)(593));                                                         
                                                                                                                                     
        global_tmr_voter(2)(594)  <=    (tmr_registers(0)(594) and tmr_registers(1)(594)) or                                            
                            (tmr_registers(1)(594) and tmr_registers(2)(594)) or                                                       
                            (tmr_registers(0)(594) and tmr_registers(2)(594));                                                         
                                                                                                                                     
        global_tmr_voter(2)(595)  <=    (tmr_registers(0)(595) and tmr_registers(1)(595)) or                                            
                            (tmr_registers(1)(595) and tmr_registers(2)(595)) or                                                       
                            (tmr_registers(0)(595) and tmr_registers(2)(595));                                                         
                                                                                                                                     
        global_tmr_voter(2)(596)  <=    (tmr_registers(0)(596) and tmr_registers(1)(596)) or                                            
                            (tmr_registers(1)(596) and tmr_registers(2)(596)) or                                                       
                            (tmr_registers(0)(596) and tmr_registers(2)(596));                                                         
                                                                                                                                     
        global_tmr_voter(2)(597)  <=    (tmr_registers(0)(597) and tmr_registers(1)(597)) or                                            
                            (tmr_registers(1)(597) and tmr_registers(2)(597)) or                                                       
                            (tmr_registers(0)(597) and tmr_registers(2)(597));                                                         
                                                                                                                                     
        global_tmr_voter(2)(598)  <=    (tmr_registers(0)(598) and tmr_registers(1)(598)) or                                            
                            (tmr_registers(1)(598) and tmr_registers(2)(598)) or                                                       
                            (tmr_registers(0)(598) and tmr_registers(2)(598));                                                         
                                                                                                                                     
        global_tmr_voter(2)(599)  <=    (tmr_registers(0)(599) and tmr_registers(1)(599)) or                                            
                            (tmr_registers(1)(599) and tmr_registers(2)(599)) or                                                       
                            (tmr_registers(0)(599) and tmr_registers(2)(599));                                                         
                                                                                                                                     
        global_tmr_voter(2)(600)  <=    (tmr_registers(0)(600) and tmr_registers(1)(600)) or                                            
                            (tmr_registers(1)(600) and tmr_registers(2)(600)) or                                                       
                            (tmr_registers(0)(600) and tmr_registers(2)(600));                                                         
                                                                                                                                     
        global_tmr_voter(2)(601)  <=    (tmr_registers(0)(601) and tmr_registers(1)(601)) or                                            
                            (tmr_registers(1)(601) and tmr_registers(2)(601)) or                                                       
                            (tmr_registers(0)(601) and tmr_registers(2)(601));                                                         
                                                                                                                                     
        global_tmr_voter(2)(602)  <=    (tmr_registers(0)(602) and tmr_registers(1)(602)) or                                            
                            (tmr_registers(1)(602) and tmr_registers(2)(602)) or                                                       
                            (tmr_registers(0)(602) and tmr_registers(2)(602));                                                         
                                                                                                                                     
        global_tmr_voter(2)(603)  <=    (tmr_registers(0)(603) and tmr_registers(1)(603)) or                                            
                            (tmr_registers(1)(603) and tmr_registers(2)(603)) or                                                       
                            (tmr_registers(0)(603) and tmr_registers(2)(603));                                                         
                                                                                                                                     
        global_tmr_voter(2)(604)  <=    (tmr_registers(0)(604) and tmr_registers(1)(604)) or                                            
                            (tmr_registers(1)(604) and tmr_registers(2)(604)) or                                                       
                            (tmr_registers(0)(604) and tmr_registers(2)(604));                                                         
                                                                                                                                     
        global_tmr_voter(2)(605)  <=    (tmr_registers(0)(605) and tmr_registers(1)(605)) or                                            
                            (tmr_registers(1)(605) and tmr_registers(2)(605)) or                                                       
                            (tmr_registers(0)(605) and tmr_registers(2)(605));                                                         
                                                                                                                                     
        global_tmr_voter(2)(606)  <=    (tmr_registers(0)(606) and tmr_registers(1)(606)) or                                            
                            (tmr_registers(1)(606) and tmr_registers(2)(606)) or                                                       
                            (tmr_registers(0)(606) and tmr_registers(2)(606));                                                         
                                                                                                                                     
        global_tmr_voter(2)(607)  <=    (tmr_registers(0)(607) and tmr_registers(1)(607)) or                                            
                            (tmr_registers(1)(607) and tmr_registers(2)(607)) or                                                       
                            (tmr_registers(0)(607) and tmr_registers(2)(607));                                                         
                                                                                                                                     
        global_tmr_voter(2)(608)  <=    (tmr_registers(0)(608) and tmr_registers(1)(608)) or                                            
                            (tmr_registers(1)(608) and tmr_registers(2)(608)) or                                                       
                            (tmr_registers(0)(608) and tmr_registers(2)(608));                                                         
                                                                                                                                     
        global_tmr_voter(2)(609)  <=    (tmr_registers(0)(609) and tmr_registers(1)(609)) or                                            
                            (tmr_registers(1)(609) and tmr_registers(2)(609)) or                                                       
                            (tmr_registers(0)(609) and tmr_registers(2)(609));                                                         
                                                                                                                                     
        global_tmr_voter(2)(610)  <=    (tmr_registers(0)(610) and tmr_registers(1)(610)) or                                            
                            (tmr_registers(1)(610) and tmr_registers(2)(610)) or                                                       
                            (tmr_registers(0)(610) and tmr_registers(2)(610));                                                         
                                                                                                                                     
        global_tmr_voter(2)(611)  <=    (tmr_registers(0)(611) and tmr_registers(1)(611)) or                                            
                            (tmr_registers(1)(611) and tmr_registers(2)(611)) or                                                       
                            (tmr_registers(0)(611) and tmr_registers(2)(611));                                                         
                                                                                                                                     
        global_tmr_voter(2)(612)  <=    (tmr_registers(0)(612) and tmr_registers(1)(612)) or                                            
                            (tmr_registers(1)(612) and tmr_registers(2)(612)) or                                                       
                            (tmr_registers(0)(612) and tmr_registers(2)(612));                                                         
                                                                                                                                     
        global_tmr_voter(2)(613)  <=    (tmr_registers(0)(613) and tmr_registers(1)(613)) or                                            
                            (tmr_registers(1)(613) and tmr_registers(2)(613)) or                                                       
                            (tmr_registers(0)(613) and tmr_registers(2)(613));                                                         
                                                                                                                                     
        global_tmr_voter(2)(614)  <=    (tmr_registers(0)(614) and tmr_registers(1)(614)) or                                            
                            (tmr_registers(1)(614) and tmr_registers(2)(614)) or                                                       
                            (tmr_registers(0)(614) and tmr_registers(2)(614));                                                         
                                                                                                                                     
        global_tmr_voter(2)(615)  <=    (tmr_registers(0)(615) and tmr_registers(1)(615)) or                                            
                            (tmr_registers(1)(615) and tmr_registers(2)(615)) or                                                       
                            (tmr_registers(0)(615) and tmr_registers(2)(615));                                                         
                                                                                                                                     
        global_tmr_voter(2)(616)  <=    (tmr_registers(0)(616) and tmr_registers(1)(616)) or                                            
                            (tmr_registers(1)(616) and tmr_registers(2)(616)) or                                                       
                            (tmr_registers(0)(616) and tmr_registers(2)(616));                                                         
                                                                                                                                     
        global_tmr_voter(2)(617)  <=    (tmr_registers(0)(617) and tmr_registers(1)(617)) or                                            
                            (tmr_registers(1)(617) and tmr_registers(2)(617)) or                                                       
                            (tmr_registers(0)(617) and tmr_registers(2)(617));                                                         
                                                                                                                                     
        global_tmr_voter(2)(618)  <=    (tmr_registers(0)(618) and tmr_registers(1)(618)) or                                            
                            (tmr_registers(1)(618) and tmr_registers(2)(618)) or                                                       
                            (tmr_registers(0)(618) and tmr_registers(2)(618));                                                         
                                                                                                                                     
        global_tmr_voter(2)(619)  <=    (tmr_registers(0)(619) and tmr_registers(1)(619)) or                                            
                            (tmr_registers(1)(619) and tmr_registers(2)(619)) or                                                       
                            (tmr_registers(0)(619) and tmr_registers(2)(619));                                                         
                                                                                                                                     
        global_tmr_voter(2)(620)  <=    (tmr_registers(0)(620) and tmr_registers(1)(620)) or                                            
                            (tmr_registers(1)(620) and tmr_registers(2)(620)) or                                                       
                            (tmr_registers(0)(620) and tmr_registers(2)(620));                                                         
                                                                                                                                     
        global_tmr_voter(2)(621)  <=    (tmr_registers(0)(621) and tmr_registers(1)(621)) or                                            
                            (tmr_registers(1)(621) and tmr_registers(2)(621)) or                                                       
                            (tmr_registers(0)(621) and tmr_registers(2)(621));                                                         
                                                                                                                                     
        global_tmr_voter(2)(622)  <=    (tmr_registers(0)(622) and tmr_registers(1)(622)) or                                            
                            (tmr_registers(1)(622) and tmr_registers(2)(622)) or                                                       
                            (tmr_registers(0)(622) and tmr_registers(2)(622));                                                         
                                                                                                                                     
        global_tmr_voter(2)(623)  <=    (tmr_registers(0)(623) and tmr_registers(1)(623)) or                                            
                            (tmr_registers(1)(623) and tmr_registers(2)(623)) or                                                       
                            (tmr_registers(0)(623) and tmr_registers(2)(623));                                                         
                                                                                                                                     
        global_tmr_voter(2)(624)  <=    (tmr_registers(0)(624) and tmr_registers(1)(624)) or                                            
                            (tmr_registers(1)(624) and tmr_registers(2)(624)) or                                                       
                            (tmr_registers(0)(624) and tmr_registers(2)(624));                                                         
                                                                                                                                     
        global_tmr_voter(2)(625)  <=    (tmr_registers(0)(625) and tmr_registers(1)(625)) or                                            
                            (tmr_registers(1)(625) and tmr_registers(2)(625)) or                                                       
                            (tmr_registers(0)(625) and tmr_registers(2)(625));                                                         
                                                                                                                                     
        global_tmr_voter(2)(626)  <=    (tmr_registers(0)(626) and tmr_registers(1)(626)) or                                            
                            (tmr_registers(1)(626) and tmr_registers(2)(626)) or                                                       
                            (tmr_registers(0)(626) and tmr_registers(2)(626));                                                         
                                                                                                                                     
        global_tmr_voter(2)(627)  <=    (tmr_registers(0)(627) and tmr_registers(1)(627)) or                                            
                            (tmr_registers(1)(627) and tmr_registers(2)(627)) or                                                       
                            (tmr_registers(0)(627) and tmr_registers(2)(627));                                                         
                                                                                                                                     
        global_tmr_voter(2)(628)  <=    (tmr_registers(0)(628) and tmr_registers(1)(628)) or                                            
                            (tmr_registers(1)(628) and tmr_registers(2)(628)) or                                                       
                            (tmr_registers(0)(628) and tmr_registers(2)(628));                                                         
                                                                                                                                     
        global_tmr_voter(2)(629)  <=    (tmr_registers(0)(629) and tmr_registers(1)(629)) or                                            
                            (tmr_registers(1)(629) and tmr_registers(2)(629)) or                                                       
                            (tmr_registers(0)(629) and tmr_registers(2)(629));                                                         
                                                                                                                                     
        global_tmr_voter(2)(630)  <=    (tmr_registers(0)(630) and tmr_registers(1)(630)) or                                            
                            (tmr_registers(1)(630) and tmr_registers(2)(630)) or                                                       
                            (tmr_registers(0)(630) and tmr_registers(2)(630));                                                         
                                                                                                                                     
        global_tmr_voter(2)(631)  <=    (tmr_registers(0)(631) and tmr_registers(1)(631)) or                                            
                            (tmr_registers(1)(631) and tmr_registers(2)(631)) or                                                       
                            (tmr_registers(0)(631) and tmr_registers(2)(631));                                                         
                                                                                                                                     
        global_tmr_voter(2)(632)  <=    (tmr_registers(0)(632) and tmr_registers(1)(632)) or                                            
                            (tmr_registers(1)(632) and tmr_registers(2)(632)) or                                                       
                            (tmr_registers(0)(632) and tmr_registers(2)(632));                                                         
                                                                                                                                     
        global_tmr_voter(2)(633)  <=    (tmr_registers(0)(633) and tmr_registers(1)(633)) or                                            
                            (tmr_registers(1)(633) and tmr_registers(2)(633)) or                                                       
                            (tmr_registers(0)(633) and tmr_registers(2)(633));                                                         
                                                                                                                                     
        global_tmr_voter(2)(634)  <=    (tmr_registers(0)(634) and tmr_registers(1)(634)) or                                            
                            (tmr_registers(1)(634) and tmr_registers(2)(634)) or                                                       
                            (tmr_registers(0)(634) and tmr_registers(2)(634));                                                         
                                                                                                                                     
        global_tmr_voter(2)(635)  <=    (tmr_registers(0)(635) and tmr_registers(1)(635)) or                                            
                            (tmr_registers(1)(635) and tmr_registers(2)(635)) or                                                       
                            (tmr_registers(0)(635) and tmr_registers(2)(635));                                                         
                                                                                                                                     
        global_tmr_voter(2)(636)  <=    (tmr_registers(0)(636) and tmr_registers(1)(636)) or                                            
                            (tmr_registers(1)(636) and tmr_registers(2)(636)) or                                                       
                            (tmr_registers(0)(636) and tmr_registers(2)(636));                                                         
                                                                                                                                     
        global_tmr_voter(2)(637)  <=    (tmr_registers(0)(637) and tmr_registers(1)(637)) or                                            
                            (tmr_registers(1)(637) and tmr_registers(2)(637)) or                                                       
                            (tmr_registers(0)(637) and tmr_registers(2)(637));                                                         
                                                                                                                                     
        global_tmr_voter(2)(638)  <=    (tmr_registers(0)(638) and tmr_registers(1)(638)) or                                            
                            (tmr_registers(1)(638) and tmr_registers(2)(638)) or                                                       
                            (tmr_registers(0)(638) and tmr_registers(2)(638));                                                         
                                                                                                                                     
        global_tmr_voter(2)(639)  <=    (tmr_registers(0)(639) and tmr_registers(1)(639)) or                                            
                            (tmr_registers(1)(639) and tmr_registers(2)(639)) or                                                       
                            (tmr_registers(0)(639) and tmr_registers(2)(639));                                                         
                                                                                                                                     
        global_tmr_voter(2)(640)  <=    (tmr_registers(0)(640) and tmr_registers(1)(640)) or                                            
                            (tmr_registers(1)(640) and tmr_registers(2)(640)) or                                                       
                            (tmr_registers(0)(640) and tmr_registers(2)(640));                                                         
                                                                                                                                     
        global_tmr_voter(2)(641)  <=    (tmr_registers(0)(641) and tmr_registers(1)(641)) or                                            
                            (tmr_registers(1)(641) and tmr_registers(2)(641)) or                                                       
                            (tmr_registers(0)(641) and tmr_registers(2)(641));                                                         
                                                                                                                                     
        global_tmr_voter(2)(642)  <=    (tmr_registers(0)(642) and tmr_registers(1)(642)) or                                            
                            (tmr_registers(1)(642) and tmr_registers(2)(642)) or                                                       
                            (tmr_registers(0)(642) and tmr_registers(2)(642));                                                         
                                                                                                                                     
        global_tmr_voter(2)(643)  <=    (tmr_registers(0)(643) and tmr_registers(1)(643)) or                                            
                            (tmr_registers(1)(643) and tmr_registers(2)(643)) or                                                       
                            (tmr_registers(0)(643) and tmr_registers(2)(643));                                                         
                                                                                                                                     
        global_tmr_voter(2)(644)  <=    (tmr_registers(0)(644) and tmr_registers(1)(644)) or                                            
                            (tmr_registers(1)(644) and tmr_registers(2)(644)) or                                                       
                            (tmr_registers(0)(644) and tmr_registers(2)(644));                                                         
                                                                                                                                     
        global_tmr_voter(2)(645)  <=    (tmr_registers(0)(645) and tmr_registers(1)(645)) or                                            
                            (tmr_registers(1)(645) and tmr_registers(2)(645)) or                                                       
                            (tmr_registers(0)(645) and tmr_registers(2)(645));                                                         
                                                                                                                                     
        global_tmr_voter(2)(646)  <=    (tmr_registers(0)(646) and tmr_registers(1)(646)) or                                            
                            (tmr_registers(1)(646) and tmr_registers(2)(646)) or                                                       
                            (tmr_registers(0)(646) and tmr_registers(2)(646));                                                         
                                                                                                                                     
        global_tmr_voter(2)(647)  <=    (tmr_registers(0)(647) and tmr_registers(1)(647)) or                                            
                            (tmr_registers(1)(647) and tmr_registers(2)(647)) or                                                       
                            (tmr_registers(0)(647) and tmr_registers(2)(647));                                                         
                                                                                                                                     
        global_tmr_voter(2)(648)  <=    (tmr_registers(0)(648) and tmr_registers(1)(648)) or                                            
                            (tmr_registers(1)(648) and tmr_registers(2)(648)) or                                                       
                            (tmr_registers(0)(648) and tmr_registers(2)(648));                                                         
                                                                                                                                     
        global_tmr_voter(2)(649)  <=    (tmr_registers(0)(649) and tmr_registers(1)(649)) or                                            
                            (tmr_registers(1)(649) and tmr_registers(2)(649)) or                                                       
                            (tmr_registers(0)(649) and tmr_registers(2)(649));                                                         
                                                                                                                                     
        global_tmr_voter(2)(650)  <=    (tmr_registers(0)(650) and tmr_registers(1)(650)) or                                            
                            (tmr_registers(1)(650) and tmr_registers(2)(650)) or                                                       
                            (tmr_registers(0)(650) and tmr_registers(2)(650));                                                         
                                                                                                                                     
        global_tmr_voter(2)(651)  <=    (tmr_registers(0)(651) and tmr_registers(1)(651)) or                                            
                            (tmr_registers(1)(651) and tmr_registers(2)(651)) or                                                       
                            (tmr_registers(0)(651) and tmr_registers(2)(651));                                                         
                                                                                                                                     
        global_tmr_voter(2)(652)  <=    (tmr_registers(0)(652) and tmr_registers(1)(652)) or                                            
                            (tmr_registers(1)(652) and tmr_registers(2)(652)) or                                                       
                            (tmr_registers(0)(652) and tmr_registers(2)(652));                                                         
                                                                                                                                     
        global_tmr_voter(2)(653)  <=    (tmr_registers(0)(653) and tmr_registers(1)(653)) or                                            
                            (tmr_registers(1)(653) and tmr_registers(2)(653)) or                                                       
                            (tmr_registers(0)(653) and tmr_registers(2)(653));                                                         
                                                                                                                                     
        global_tmr_voter(2)(654)  <=    (tmr_registers(0)(654) and tmr_registers(1)(654)) or                                            
                            (tmr_registers(1)(654) and tmr_registers(2)(654)) or                                                       
                            (tmr_registers(0)(654) and tmr_registers(2)(654));                                                         
                                                                                                                                     
        global_tmr_voter(2)(655)  <=    (tmr_registers(0)(655) and tmr_registers(1)(655)) or                                            
                            (tmr_registers(1)(655) and tmr_registers(2)(655)) or                                                       
                            (tmr_registers(0)(655) and tmr_registers(2)(655));                                                         
                                                                                                                                     
        global_tmr_voter(2)(656)  <=    (tmr_registers(0)(656) and tmr_registers(1)(656)) or                                            
                            (tmr_registers(1)(656) and tmr_registers(2)(656)) or                                                       
                            (tmr_registers(0)(656) and tmr_registers(2)(656));                                                         
                                                                                                                                     
        global_tmr_voter(2)(657)  <=    (tmr_registers(0)(657) and tmr_registers(1)(657)) or                                            
                            (tmr_registers(1)(657) and tmr_registers(2)(657)) or                                                       
                            (tmr_registers(0)(657) and tmr_registers(2)(657));                                                         
                                                                                                                                     
        global_tmr_voter(2)(658)  <=    (tmr_registers(0)(658) and tmr_registers(1)(658)) or                                            
                            (tmr_registers(1)(658) and tmr_registers(2)(658)) or                                                       
                            (tmr_registers(0)(658) and tmr_registers(2)(658));                                                         
                                                                                                                                     
        global_tmr_voter(2)(659)  <=    (tmr_registers(0)(659) and tmr_registers(1)(659)) or                                            
                            (tmr_registers(1)(659) and tmr_registers(2)(659)) or                                                       
                            (tmr_registers(0)(659) and tmr_registers(2)(659));                                                         
                                                                                                                                     
        global_tmr_voter(2)(660)  <=    (tmr_registers(0)(660) and tmr_registers(1)(660)) or                                            
                            (tmr_registers(1)(660) and tmr_registers(2)(660)) or                                                       
                            (tmr_registers(0)(660) and tmr_registers(2)(660));                                                         
                                                                                                                                     
        global_tmr_voter(2)(661)  <=    (tmr_registers(0)(661) and tmr_registers(1)(661)) or                                            
                            (tmr_registers(1)(661) and tmr_registers(2)(661)) or                                                       
                            (tmr_registers(0)(661) and tmr_registers(2)(661));                                                         
                                                                                                                                     
        global_tmr_voter(2)(662)  <=    (tmr_registers(0)(662) and tmr_registers(1)(662)) or                                            
                            (tmr_registers(1)(662) and tmr_registers(2)(662)) or                                                       
                            (tmr_registers(0)(662) and tmr_registers(2)(662));                                                         
                                                                                                                                     
        global_tmr_voter(2)(663)  <=    (tmr_registers(0)(663) and tmr_registers(1)(663)) or                                            
                            (tmr_registers(1)(663) and tmr_registers(2)(663)) or                                                       
                            (tmr_registers(0)(663) and tmr_registers(2)(663));                                                         
                                                                                                                                     
        global_tmr_voter(2)(664)  <=    (tmr_registers(0)(664) and tmr_registers(1)(664)) or                                            
                            (tmr_registers(1)(664) and tmr_registers(2)(664)) or                                                       
                            (tmr_registers(0)(664) and tmr_registers(2)(664));                                                         
                                                                                                                                     
        global_tmr_voter(2)(665)  <=    (tmr_registers(0)(665) and tmr_registers(1)(665)) or                                            
                            (tmr_registers(1)(665) and tmr_registers(2)(665)) or                                                       
                            (tmr_registers(0)(665) and tmr_registers(2)(665));                                                         
                                                                                                                                     
        global_tmr_voter(2)(666)  <=    (tmr_registers(0)(666) and tmr_registers(1)(666)) or                                            
                            (tmr_registers(1)(666) and tmr_registers(2)(666)) or                                                       
                            (tmr_registers(0)(666) and tmr_registers(2)(666));                                                         
                                                                                                                                     
        global_tmr_voter(2)(667)  <=    (tmr_registers(0)(667) and tmr_registers(1)(667)) or                                            
                            (tmr_registers(1)(667) and tmr_registers(2)(667)) or                                                       
                            (tmr_registers(0)(667) and tmr_registers(2)(667));                                                         
                                                                                                                                     
        global_tmr_voter(2)(668)  <=    (tmr_registers(0)(668) and tmr_registers(1)(668)) or                                            
                            (tmr_registers(1)(668) and tmr_registers(2)(668)) or                                                       
                            (tmr_registers(0)(668) and tmr_registers(2)(668));                                                         
                                                                                                                                     
        global_tmr_voter(2)(669)  <=    (tmr_registers(0)(669) and tmr_registers(1)(669)) or                                            
                            (tmr_registers(1)(669) and tmr_registers(2)(669)) or                                                       
                            (tmr_registers(0)(669) and tmr_registers(2)(669));                                                         
                                                                                                                                     
        global_tmr_voter(2)(670)  <=    (tmr_registers(0)(670) and tmr_registers(1)(670)) or                                            
                            (tmr_registers(1)(670) and tmr_registers(2)(670)) or                                                       
                            (tmr_registers(0)(670) and tmr_registers(2)(670));                                                         
                                                                                                                                     
        global_tmr_voter(2)(671)  <=    (tmr_registers(0)(671) and tmr_registers(1)(671)) or                                            
                            (tmr_registers(1)(671) and tmr_registers(2)(671)) or                                                       
                            (tmr_registers(0)(671) and tmr_registers(2)(671));                                                         
                                                                                                                                     
        global_tmr_voter(2)(672)  <=    (tmr_registers(0)(672) and tmr_registers(1)(672)) or                                            
                            (tmr_registers(1)(672) and tmr_registers(2)(672)) or                                                       
                            (tmr_registers(0)(672) and tmr_registers(2)(672));                                                         
                                                                                                                                     
        global_tmr_voter(2)(673)  <=    (tmr_registers(0)(673) and tmr_registers(1)(673)) or                                            
                            (tmr_registers(1)(673) and tmr_registers(2)(673)) or                                                       
                            (tmr_registers(0)(673) and tmr_registers(2)(673));                                                         
                                                                                                                                     
        global_tmr_voter(2)(674)  <=    (tmr_registers(0)(674) and tmr_registers(1)(674)) or                                            
                            (tmr_registers(1)(674) and tmr_registers(2)(674)) or                                                       
                            (tmr_registers(0)(674) and tmr_registers(2)(674));                                                         
                                                                                                                                     
        global_tmr_voter(2)(675)  <=    (tmr_registers(0)(675) and tmr_registers(1)(675)) or                                            
                            (tmr_registers(1)(675) and tmr_registers(2)(675)) or                                                       
                            (tmr_registers(0)(675) and tmr_registers(2)(675));                                                         
                                                                                                                                     
        global_tmr_voter(2)(676)  <=    (tmr_registers(0)(676) and tmr_registers(1)(676)) or                                            
                            (tmr_registers(1)(676) and tmr_registers(2)(676)) or                                                       
                            (tmr_registers(0)(676) and tmr_registers(2)(676));                                                         
                                                                                                                                     
        global_tmr_voter(2)(677)  <=    (tmr_registers(0)(677) and tmr_registers(1)(677)) or                                            
                            (tmr_registers(1)(677) and tmr_registers(2)(677)) or                                                       
                            (tmr_registers(0)(677) and tmr_registers(2)(677));                                                         
                                                                                                                                     
        global_tmr_voter(2)(678)  <=    (tmr_registers(0)(678) and tmr_registers(1)(678)) or                                            
                            (tmr_registers(1)(678) and tmr_registers(2)(678)) or                                                       
                            (tmr_registers(0)(678) and tmr_registers(2)(678));                                                         
                                                                                                                                     
        global_tmr_voter(2)(679)  <=    (tmr_registers(0)(679) and tmr_registers(1)(679)) or                                            
                            (tmr_registers(1)(679) and tmr_registers(2)(679)) or                                                       
                            (tmr_registers(0)(679) and tmr_registers(2)(679));                                                         
                                                                                                                                     
        global_tmr_voter(2)(680)  <=    (tmr_registers(0)(680) and tmr_registers(1)(680)) or                                            
                            (tmr_registers(1)(680) and tmr_registers(2)(680)) or                                                       
                            (tmr_registers(0)(680) and tmr_registers(2)(680));                                                         
                                                                                                                                     
        global_tmr_voter(2)(681)  <=    (tmr_registers(0)(681) and tmr_registers(1)(681)) or                                            
                            (tmr_registers(1)(681) and tmr_registers(2)(681)) or                                                       
                            (tmr_registers(0)(681) and tmr_registers(2)(681));                                                         
                                                                                                                                     
        global_tmr_voter(2)(682)  <=    (tmr_registers(0)(682) and tmr_registers(1)(682)) or                                            
                            (tmr_registers(1)(682) and tmr_registers(2)(682)) or                                                       
                            (tmr_registers(0)(682) and tmr_registers(2)(682));                                                         
                                                                                                                                     
        global_tmr_voter(2)(683)  <=    (tmr_registers(0)(683) and tmr_registers(1)(683)) or                                            
                            (tmr_registers(1)(683) and tmr_registers(2)(683)) or                                                       
                            (tmr_registers(0)(683) and tmr_registers(2)(683));                                                         
                                                                                                                                     
        global_tmr_voter(2)(684)  <=    (tmr_registers(0)(684) and tmr_registers(1)(684)) or                                            
                            (tmr_registers(1)(684) and tmr_registers(2)(684)) or                                                       
                            (tmr_registers(0)(684) and tmr_registers(2)(684));                                                         
                                                                                                                                     
        global_tmr_voter(2)(685)  <=    (tmr_registers(0)(685) and tmr_registers(1)(685)) or                                            
                            (tmr_registers(1)(685) and tmr_registers(2)(685)) or                                                       
                            (tmr_registers(0)(685) and tmr_registers(2)(685));                                                         
                                                                                                                                     
        global_tmr_voter(2)(686)  <=    (tmr_registers(0)(686) and tmr_registers(1)(686)) or                                            
                            (tmr_registers(1)(686) and tmr_registers(2)(686)) or                                                       
                            (tmr_registers(0)(686) and tmr_registers(2)(686));                                                         
                                                                                                                                     
        global_tmr_voter(2)(687)  <=    (tmr_registers(0)(687) and tmr_registers(1)(687)) or                                            
                            (tmr_registers(1)(687) and tmr_registers(2)(687)) or                                                       
                            (tmr_registers(0)(687) and tmr_registers(2)(687));                                                         
                                                                                                                                     
        global_tmr_voter(2)(688)  <=    (tmr_registers(0)(688) and tmr_registers(1)(688)) or                                            
                            (tmr_registers(1)(688) and tmr_registers(2)(688)) or                                                       
                            (tmr_registers(0)(688) and tmr_registers(2)(688));                                                         
                                                                                                                                     
        global_tmr_voter(2)(689)  <=    (tmr_registers(0)(689) and tmr_registers(1)(689)) or                                            
                            (tmr_registers(1)(689) and tmr_registers(2)(689)) or                                                       
                            (tmr_registers(0)(689) and tmr_registers(2)(689));                                                         
                                                                                                                                     
        global_tmr_voter(2)(690)  <=    (tmr_registers(0)(690) and tmr_registers(1)(690)) or                                            
                            (tmr_registers(1)(690) and tmr_registers(2)(690)) or                                                       
                            (tmr_registers(0)(690) and tmr_registers(2)(690));                                                         
                                                                                                                                     
        global_tmr_voter(2)(691)  <=    (tmr_registers(0)(691) and tmr_registers(1)(691)) or                                            
                            (tmr_registers(1)(691) and tmr_registers(2)(691)) or                                                       
                            (tmr_registers(0)(691) and tmr_registers(2)(691));                                                         
                                                                                                                                     
        global_tmr_voter(2)(692)  <=    (tmr_registers(0)(692) and tmr_registers(1)(692)) or                                            
                            (tmr_registers(1)(692) and tmr_registers(2)(692)) or                                                       
                            (tmr_registers(0)(692) and tmr_registers(2)(692));                                                         
                                                                                                                                     
        global_tmr_voter(2)(693)  <=    (tmr_registers(0)(693) and tmr_registers(1)(693)) or                                            
                            (tmr_registers(1)(693) and tmr_registers(2)(693)) or                                                       
                            (tmr_registers(0)(693) and tmr_registers(2)(693));                                                         
                                                                                                                                     
        global_tmr_voter(2)(694)  <=    (tmr_registers(0)(694) and tmr_registers(1)(694)) or                                            
                            (tmr_registers(1)(694) and tmr_registers(2)(694)) or                                                       
                            (tmr_registers(0)(694) and tmr_registers(2)(694));                                                         
                                                                                                                                     
        global_tmr_voter(2)(695)  <=    (tmr_registers(0)(695) and tmr_registers(1)(695)) or                                            
                            (tmr_registers(1)(695) and tmr_registers(2)(695)) or                                                       
                            (tmr_registers(0)(695) and tmr_registers(2)(695));                                                         
                                                                                                                                     
        global_tmr_voter(2)(696)  <=    (tmr_registers(0)(696) and tmr_registers(1)(696)) or                                            
                            (tmr_registers(1)(696) and tmr_registers(2)(696)) or                                                       
                            (tmr_registers(0)(696) and tmr_registers(2)(696));                                                         
                                                                                                                                     
        global_tmr_voter(2)(697)  <=    (tmr_registers(0)(697) and tmr_registers(1)(697)) or                                            
                            (tmr_registers(1)(697) and tmr_registers(2)(697)) or                                                       
                            (tmr_registers(0)(697) and tmr_registers(2)(697));                                                         
                                                                                                                                     
        global_tmr_voter(2)(698)  <=    (tmr_registers(0)(698) and tmr_registers(1)(698)) or                                            
                            (tmr_registers(1)(698) and tmr_registers(2)(698)) or                                                       
                            (tmr_registers(0)(698) and tmr_registers(2)(698));                                                         
                                                                                                                                     
        global_tmr_voter(2)(699)  <=    (tmr_registers(0)(699) and tmr_registers(1)(699)) or                                            
                            (tmr_registers(1)(699) and tmr_registers(2)(699)) or                                                       
                            (tmr_registers(0)(699) and tmr_registers(2)(699));                                                         
                                                                                                                                     
        global_tmr_voter(2)(700)  <=    (tmr_registers(0)(700) and tmr_registers(1)(700)) or                                            
                            (tmr_registers(1)(700) and tmr_registers(2)(700)) or                                                       
                            (tmr_registers(0)(700) and tmr_registers(2)(700));                                                         
                                                                                                                                     
        global_tmr_voter(2)(701)  <=    (tmr_registers(0)(701) and tmr_registers(1)(701)) or                                            
                            (tmr_registers(1)(701) and tmr_registers(2)(701)) or                                                       
                            (tmr_registers(0)(701) and tmr_registers(2)(701));                                                         
                                                                                                                                     
        global_tmr_voter(2)(702)  <=    (tmr_registers(0)(702) and tmr_registers(1)(702)) or                                            
                            (tmr_registers(1)(702) and tmr_registers(2)(702)) or                                                       
                            (tmr_registers(0)(702) and tmr_registers(2)(702));                                                         
                                                                                                                                     
        global_tmr_voter(2)(703)  <=    (tmr_registers(0)(703) and tmr_registers(1)(703)) or                                            
                            (tmr_registers(1)(703) and tmr_registers(2)(703)) or                                                       
                            (tmr_registers(0)(703) and tmr_registers(2)(703));                                                         
                                                                                                                                     
        global_tmr_voter(2)(704)  <=    (tmr_registers(0)(704) and tmr_registers(1)(704)) or                                            
                            (tmr_registers(1)(704) and tmr_registers(2)(704)) or                                                       
                            (tmr_registers(0)(704) and tmr_registers(2)(704));                                                         
                                                                                                                                     
        global_tmr_voter(2)(705)  <=    (tmr_registers(0)(705) and tmr_registers(1)(705)) or                                            
                            (tmr_registers(1)(705) and tmr_registers(2)(705)) or                                                       
                            (tmr_registers(0)(705) and tmr_registers(2)(705));                                                         
                                                                                                                                     
        global_tmr_voter(2)(706)  <=    (tmr_registers(0)(706) and tmr_registers(1)(706)) or                                            
                            (tmr_registers(1)(706) and tmr_registers(2)(706)) or                                                       
                            (tmr_registers(0)(706) and tmr_registers(2)(706));                                                         
                                                                                                                                     
        global_tmr_voter(2)(707)  <=    (tmr_registers(0)(707) and tmr_registers(1)(707)) or                                            
                            (tmr_registers(1)(707) and tmr_registers(2)(707)) or                                                       
                            (tmr_registers(0)(707) and tmr_registers(2)(707));                                                         
                                                                                                                                     
        global_tmr_voter(2)(708)  <=    (tmr_registers(0)(708) and tmr_registers(1)(708)) or                                            
                            (tmr_registers(1)(708) and tmr_registers(2)(708)) or                                                       
                            (tmr_registers(0)(708) and tmr_registers(2)(708));                                                         
                                                                                                                                     
        global_tmr_voter(2)(709)  <=    (tmr_registers(0)(709) and tmr_registers(1)(709)) or                                            
                            (tmr_registers(1)(709) and tmr_registers(2)(709)) or                                                       
                            (tmr_registers(0)(709) and tmr_registers(2)(709));                                                         
                                                                                                                                     
        global_tmr_voter(2)(710)  <=    (tmr_registers(0)(710) and tmr_registers(1)(710)) or                                            
                            (tmr_registers(1)(710) and tmr_registers(2)(710)) or                                                       
                            (tmr_registers(0)(710) and tmr_registers(2)(710));                                                         
                                                                                                                                     
        global_tmr_voter(2)(711)  <=    (tmr_registers(0)(711) and tmr_registers(1)(711)) or                                            
                            (tmr_registers(1)(711) and tmr_registers(2)(711)) or                                                       
                            (tmr_registers(0)(711) and tmr_registers(2)(711));                                                         
                                                                                                                                     
        global_tmr_voter(2)(712)  <=    (tmr_registers(0)(712) and tmr_registers(1)(712)) or                                            
                            (tmr_registers(1)(712) and tmr_registers(2)(712)) or                                                       
                            (tmr_registers(0)(712) and tmr_registers(2)(712));                                                         
                                                                                                                                     
        global_tmr_voter(2)(713)  <=    (tmr_registers(0)(713) and tmr_registers(1)(713)) or                                            
                            (tmr_registers(1)(713) and tmr_registers(2)(713)) or                                                       
                            (tmr_registers(0)(713) and tmr_registers(2)(713));                                                         
                                                                                                                                     
        global_tmr_voter(2)(714)  <=    (tmr_registers(0)(714) and tmr_registers(1)(714)) or                                            
                            (tmr_registers(1)(714) and tmr_registers(2)(714)) or                                                       
                            (tmr_registers(0)(714) and tmr_registers(2)(714));                                                         
                                                                                                                                     
        global_tmr_voter(2)(715)  <=    (tmr_registers(0)(715) and tmr_registers(1)(715)) or                                            
                            (tmr_registers(1)(715) and tmr_registers(2)(715)) or                                                       
                            (tmr_registers(0)(715) and tmr_registers(2)(715));                                                         
                                                                                                                                     
        global_tmr_voter(2)(716)  <=    (tmr_registers(0)(716) and tmr_registers(1)(716)) or                                            
                            (tmr_registers(1)(716) and tmr_registers(2)(716)) or                                                       
                            (tmr_registers(0)(716) and tmr_registers(2)(716));                                                         
                                                                                                                                     
        global_tmr_voter(2)(717)  <=    (tmr_registers(0)(717) and tmr_registers(1)(717)) or                                            
                            (tmr_registers(1)(717) and tmr_registers(2)(717)) or                                                       
                            (tmr_registers(0)(717) and tmr_registers(2)(717));                                                         
                                                                                                                                     
        global_tmr_voter(2)(718)  <=    (tmr_registers(0)(718) and tmr_registers(1)(718)) or                                            
                            (tmr_registers(1)(718) and tmr_registers(2)(718)) or                                                       
                            (tmr_registers(0)(718) and tmr_registers(2)(718));                                                         
                                                                                                                                     
        global_tmr_voter(2)(719)  <=    (tmr_registers(0)(719) and tmr_registers(1)(719)) or                                            
                            (tmr_registers(1)(719) and tmr_registers(2)(719)) or                                                       
                            (tmr_registers(0)(719) and tmr_registers(2)(719));                                                         
                                                                                                                                     
        global_tmr_voter(2)(720)  <=    (tmr_registers(0)(720) and tmr_registers(1)(720)) or                                            
                            (tmr_registers(1)(720) and tmr_registers(2)(720)) or                                                       
                            (tmr_registers(0)(720) and tmr_registers(2)(720));                                                         
                                                                                                                                     
        global_tmr_voter(2)(721)  <=    (tmr_registers(0)(721) and tmr_registers(1)(721)) or                                            
                            (tmr_registers(1)(721) and tmr_registers(2)(721)) or                                                       
                            (tmr_registers(0)(721) and tmr_registers(2)(721));                                                         
                                                                                                                                     
        global_tmr_voter(2)(722)  <=    (tmr_registers(0)(722) and tmr_registers(1)(722)) or                                            
                            (tmr_registers(1)(722) and tmr_registers(2)(722)) or                                                       
                            (tmr_registers(0)(722) and tmr_registers(2)(722));                                                         
                                                                                                                                     
        global_tmr_voter(2)(723)  <=    (tmr_registers(0)(723) and tmr_registers(1)(723)) or                                            
                            (tmr_registers(1)(723) and tmr_registers(2)(723)) or                                                       
                            (tmr_registers(0)(723) and tmr_registers(2)(723));                                                         
                                                                                                                                     
        global_tmr_voter(2)(724)  <=    (tmr_registers(0)(724) and tmr_registers(1)(724)) or                                            
                            (tmr_registers(1)(724) and tmr_registers(2)(724)) or                                                       
                            (tmr_registers(0)(724) and tmr_registers(2)(724));                                                         
                                                                                                                                     
        global_tmr_voter(2)(725)  <=    (tmr_registers(0)(725) and tmr_registers(1)(725)) or                                            
                            (tmr_registers(1)(725) and tmr_registers(2)(725)) or                                                       
                            (tmr_registers(0)(725) and tmr_registers(2)(725));                                                         
                                                                                                                                     
        global_tmr_voter(2)(726)  <=    (tmr_registers(0)(726) and tmr_registers(1)(726)) or                                            
                            (tmr_registers(1)(726) and tmr_registers(2)(726)) or                                                       
                            (tmr_registers(0)(726) and tmr_registers(2)(726));                                                         
                                                                                                                                     
        global_tmr_voter(2)(727)  <=    (tmr_registers(0)(727) and tmr_registers(1)(727)) or                                            
                            (tmr_registers(1)(727) and tmr_registers(2)(727)) or                                                       
                            (tmr_registers(0)(727) and tmr_registers(2)(727));                                                         
                                                                                                                                     
        global_tmr_voter(2)(728)  <=    (tmr_registers(0)(728) and tmr_registers(1)(728)) or                                            
                            (tmr_registers(1)(728) and tmr_registers(2)(728)) or                                                       
                            (tmr_registers(0)(728) and tmr_registers(2)(728));                                                         
                                                                                                                                     
        global_tmr_voter(2)(729)  <=    (tmr_registers(0)(729) and tmr_registers(1)(729)) or                                            
                            (tmr_registers(1)(729) and tmr_registers(2)(729)) or                                                       
                            (tmr_registers(0)(729) and tmr_registers(2)(729));                                                         
                                                                                                                                     
        global_tmr_voter(2)(730)  <=    (tmr_registers(0)(730) and tmr_registers(1)(730)) or                                            
                            (tmr_registers(1)(730) and tmr_registers(2)(730)) or                                                       
                            (tmr_registers(0)(730) and tmr_registers(2)(730));                                                         
                                                                                                                                     
        global_tmr_voter(2)(731)  <=    (tmr_registers(0)(731) and tmr_registers(1)(731)) or                                            
                            (tmr_registers(1)(731) and tmr_registers(2)(731)) or                                                       
                            (tmr_registers(0)(731) and tmr_registers(2)(731));                                                         
                                                                                                                                     
        global_tmr_voter(2)(732)  <=    (tmr_registers(0)(732) and tmr_registers(1)(732)) or                                            
                            (tmr_registers(1)(732) and tmr_registers(2)(732)) or                                                       
                            (tmr_registers(0)(732) and tmr_registers(2)(732));                                                         
                                                                                                                                     
        global_tmr_voter(2)(733)  <=    (tmr_registers(0)(733) and tmr_registers(1)(733)) or                                            
                            (tmr_registers(1)(733) and tmr_registers(2)(733)) or                                                       
                            (tmr_registers(0)(733) and tmr_registers(2)(733));                                                         
                                                                                                                                     
        global_tmr_voter(2)(734)  <=    (tmr_registers(0)(734) and tmr_registers(1)(734)) or                                            
                            (tmr_registers(1)(734) and tmr_registers(2)(734)) or                                                       
                            (tmr_registers(0)(734) and tmr_registers(2)(734));                                                         
                                                                                                                                     
        global_tmr_voter(2)(735)  <=    (tmr_registers(0)(735) and tmr_registers(1)(735)) or                                            
                            (tmr_registers(1)(735) and tmr_registers(2)(735)) or                                                       
                            (tmr_registers(0)(735) and tmr_registers(2)(735));                                                         
                                                                                                                                     
        global_tmr_voter(2)(736)  <=    (tmr_registers(0)(736) and tmr_registers(1)(736)) or                                            
                            (tmr_registers(1)(736) and tmr_registers(2)(736)) or                                                       
                            (tmr_registers(0)(736) and tmr_registers(2)(736));                                                         
                                                                                                                                     
        global_tmr_voter(2)(737)  <=    (tmr_registers(0)(737) and tmr_registers(1)(737)) or                                            
                            (tmr_registers(1)(737) and tmr_registers(2)(737)) or                                                       
                            (tmr_registers(0)(737) and tmr_registers(2)(737));                                                         
                                                                                                                                     
        global_tmr_voter(2)(738)  <=    (tmr_registers(0)(738) and tmr_registers(1)(738)) or                                            
                            (tmr_registers(1)(738) and tmr_registers(2)(738)) or                                                       
                            (tmr_registers(0)(738) and tmr_registers(2)(738));                                                         
                                                                                                                                     
        global_tmr_voter(2)(739)  <=    (tmr_registers(0)(739) and tmr_registers(1)(739)) or                                            
                            (tmr_registers(1)(739) and tmr_registers(2)(739)) or                                                       
                            (tmr_registers(0)(739) and tmr_registers(2)(739));                                                         
                                                                                                                                     
        global_tmr_voter(2)(740)  <=    (tmr_registers(0)(740) and tmr_registers(1)(740)) or                                            
                            (tmr_registers(1)(740) and tmr_registers(2)(740)) or                                                       
                            (tmr_registers(0)(740) and tmr_registers(2)(740));                                                         
                                                                                                                                     
        global_tmr_voter(2)(741)  <=    (tmr_registers(0)(741) and tmr_registers(1)(741)) or                                            
                            (tmr_registers(1)(741) and tmr_registers(2)(741)) or                                                       
                            (tmr_registers(0)(741) and tmr_registers(2)(741));                                                         
                                                                                                                                     
        global_tmr_voter(2)(742)  <=    (tmr_registers(0)(742) and tmr_registers(1)(742)) or                                            
                            (tmr_registers(1)(742) and tmr_registers(2)(742)) or                                                       
                            (tmr_registers(0)(742) and tmr_registers(2)(742));                                                         
                                                                                                                                     
        global_tmr_voter(2)(743)  <=    (tmr_registers(0)(743) and tmr_registers(1)(743)) or                                            
                            (tmr_registers(1)(743) and tmr_registers(2)(743)) or                                                       
                            (tmr_registers(0)(743) and tmr_registers(2)(743));                                                         
                                                                                                                                     
        global_tmr_voter(2)(744)  <=    (tmr_registers(0)(744) and tmr_registers(1)(744)) or                                            
                            (tmr_registers(1)(744) and tmr_registers(2)(744)) or                                                       
                            (tmr_registers(0)(744) and tmr_registers(2)(744));                                                         
                                                                                                                                     
        global_tmr_voter(2)(745)  <=    (tmr_registers(0)(745) and tmr_registers(1)(745)) or                                            
                            (tmr_registers(1)(745) and tmr_registers(2)(745)) or                                                       
                            (tmr_registers(0)(745) and tmr_registers(2)(745));                                                         
                                                                                                                                     
        global_tmr_voter(2)(746)  <=    (tmr_registers(0)(746) and tmr_registers(1)(746)) or                                            
                            (tmr_registers(1)(746) and tmr_registers(2)(746)) or                                                       
                            (tmr_registers(0)(746) and tmr_registers(2)(746));                                                         
                                                                                                                                     
        global_tmr_voter(2)(747)  <=    (tmr_registers(0)(747) and tmr_registers(1)(747)) or                                            
                            (tmr_registers(1)(747) and tmr_registers(2)(747)) or                                                       
                            (tmr_registers(0)(747) and tmr_registers(2)(747));                                                         
                                                                                                                                     
        global_tmr_voter(2)(748)  <=    (tmr_registers(0)(748) and tmr_registers(1)(748)) or                                            
                            (tmr_registers(1)(748) and tmr_registers(2)(748)) or                                                       
                            (tmr_registers(0)(748) and tmr_registers(2)(748));                                                         
                                                                                                                                     
        global_tmr_voter(2)(749)  <=    (tmr_registers(0)(749) and tmr_registers(1)(749)) or                                            
                            (tmr_registers(1)(749) and tmr_registers(2)(749)) or                                                       
                            (tmr_registers(0)(749) and tmr_registers(2)(749));                                                         
                                                                                                                                     
        global_tmr_voter(2)(750)  <=    (tmr_registers(0)(750) and tmr_registers(1)(750)) or                                            
                            (tmr_registers(1)(750) and tmr_registers(2)(750)) or                                                       
                            (tmr_registers(0)(750) and tmr_registers(2)(750));                                                         
                                                                                                                                     
        global_tmr_voter(2)(751)  <=    (tmr_registers(0)(751) and tmr_registers(1)(751)) or                                            
                            (tmr_registers(1)(751) and tmr_registers(2)(751)) or                                                       
                            (tmr_registers(0)(751) and tmr_registers(2)(751));                                                         
                                                                                                                                     
        global_tmr_voter(2)(752)  <=    (tmr_registers(0)(752) and tmr_registers(1)(752)) or                                            
                            (tmr_registers(1)(752) and tmr_registers(2)(752)) or                                                       
                            (tmr_registers(0)(752) and tmr_registers(2)(752));                                                         
                                                                                                                                     
        global_tmr_voter(2)(753)  <=    (tmr_registers(0)(753) and tmr_registers(1)(753)) or                                            
                            (tmr_registers(1)(753) and tmr_registers(2)(753)) or                                                       
                            (tmr_registers(0)(753) and tmr_registers(2)(753));                                                         
                                                                                                                                     
        global_tmr_voter(2)(754)  <=    (tmr_registers(0)(754) and tmr_registers(1)(754)) or                                            
                            (tmr_registers(1)(754) and tmr_registers(2)(754)) or                                                       
                            (tmr_registers(0)(754) and tmr_registers(2)(754));                                                         
                                                                                                                                     
        global_tmr_voter(2)(755)  <=    (tmr_registers(0)(755) and tmr_registers(1)(755)) or                                            
                            (tmr_registers(1)(755) and tmr_registers(2)(755)) or                                                       
                            (tmr_registers(0)(755) and tmr_registers(2)(755));                                                         
                                                                                                                                     
        global_tmr_voter(2)(756)  <=    (tmr_registers(0)(756) and tmr_registers(1)(756)) or                                            
                            (tmr_registers(1)(756) and tmr_registers(2)(756)) or                                                       
                            (tmr_registers(0)(756) and tmr_registers(2)(756));                                                         
                                                                                                                                     
        global_tmr_voter(2)(757)  <=    (tmr_registers(0)(757) and tmr_registers(1)(757)) or                                            
                            (tmr_registers(1)(757) and tmr_registers(2)(757)) or                                                       
                            (tmr_registers(0)(757) and tmr_registers(2)(757));                                                         
                                                                                                                                     
        global_tmr_voter(2)(758)  <=    (tmr_registers(0)(758) and tmr_registers(1)(758)) or                                            
                            (tmr_registers(1)(758) and tmr_registers(2)(758)) or                                                       
                            (tmr_registers(0)(758) and tmr_registers(2)(758));                                                         
                                                                                                                                     
        global_tmr_voter(2)(759)  <=    (tmr_registers(0)(759) and tmr_registers(1)(759)) or                                            
                            (tmr_registers(1)(759) and tmr_registers(2)(759)) or                                                       
                            (tmr_registers(0)(759) and tmr_registers(2)(759));                                                         
                                                                                                                                     
        global_tmr_voter(2)(760)  <=    (tmr_registers(0)(760) and tmr_registers(1)(760)) or                                            
                            (tmr_registers(1)(760) and tmr_registers(2)(760)) or                                                       
                            (tmr_registers(0)(760) and tmr_registers(2)(760));                                                         
                                                                                                                                     
        global_tmr_voter(2)(761)  <=    (tmr_registers(0)(761) and tmr_registers(1)(761)) or                                            
                            (tmr_registers(1)(761) and tmr_registers(2)(761)) or                                                       
                            (tmr_registers(0)(761) and tmr_registers(2)(761));                                                         
                                                                                                                                     
        global_tmr_voter(2)(762)  <=    (tmr_registers(0)(762) and tmr_registers(1)(762)) or                                            
                            (tmr_registers(1)(762) and tmr_registers(2)(762)) or                                                       
                            (tmr_registers(0)(762) and tmr_registers(2)(762));                                                         
                                                                                                                                     
        global_tmr_voter(2)(763)  <=    (tmr_registers(0)(763) and tmr_registers(1)(763)) or                                            
                            (tmr_registers(1)(763) and tmr_registers(2)(763)) or                                                       
                            (tmr_registers(0)(763) and tmr_registers(2)(763));                                                         
                                                                                                                                     
        global_tmr_voter(2)(764)  <=    (tmr_registers(0)(764) and tmr_registers(1)(764)) or                                            
                            (tmr_registers(1)(764) and tmr_registers(2)(764)) or                                                       
                            (tmr_registers(0)(764) and tmr_registers(2)(764));                                                         
                                                                                                                                     
        global_tmr_voter(2)(765)  <=    (tmr_registers(0)(765) and tmr_registers(1)(765)) or                                            
                            (tmr_registers(1)(765) and tmr_registers(2)(765)) or                                                       
                            (tmr_registers(0)(765) and tmr_registers(2)(765));                                                         
                                                                                                                                     
        global_tmr_voter(2)(766)  <=    (tmr_registers(0)(766) and tmr_registers(1)(766)) or                                            
                            (tmr_registers(1)(766) and tmr_registers(2)(766)) or                                                       
                            (tmr_registers(0)(766) and tmr_registers(2)(766));                                                         
                                                                                                                                     
        global_tmr_voter(2)(767)  <=    (tmr_registers(0)(767) and tmr_registers(1)(767)) or                                            
                            (tmr_registers(1)(767) and tmr_registers(2)(767)) or                                                       
                            (tmr_registers(0)(767) and tmr_registers(2)(767));                                                         
                                                                                                                                     
        global_tmr_voter(2)(768)  <=    (tmr_registers(0)(768) and tmr_registers(1)(768)) or                                            
                            (tmr_registers(1)(768) and tmr_registers(2)(768)) or                                                       
                            (tmr_registers(0)(768) and tmr_registers(2)(768));                                                         
                                                                                                                                     
        global_tmr_voter(2)(769)  <=    (tmr_registers(0)(769) and tmr_registers(1)(769)) or                                            
                            (tmr_registers(1)(769) and tmr_registers(2)(769)) or                                                       
                            (tmr_registers(0)(769) and tmr_registers(2)(769));                                                         
                                                                                                                                     
        global_tmr_voter(2)(770)  <=    (tmr_registers(0)(770) and tmr_registers(1)(770)) or                                            
                            (tmr_registers(1)(770) and tmr_registers(2)(770)) or                                                       
                            (tmr_registers(0)(770) and tmr_registers(2)(770));                                                         
                                                                                                                                     
        global_tmr_voter(2)(771)  <=    (tmr_registers(0)(771) and tmr_registers(1)(771)) or                                            
                            (tmr_registers(1)(771) and tmr_registers(2)(771)) or                                                       
                            (tmr_registers(0)(771) and tmr_registers(2)(771));                                                         
                                                                                                                                     
        global_tmr_voter(2)(772)  <=    (tmr_registers(0)(772) and tmr_registers(1)(772)) or                                            
                            (tmr_registers(1)(772) and tmr_registers(2)(772)) or                                                       
                            (tmr_registers(0)(772) and tmr_registers(2)(772));                                                         
                                                                                                                                     
        global_tmr_voter(2)(773)  <=    (tmr_registers(0)(773) and tmr_registers(1)(773)) or                                            
                            (tmr_registers(1)(773) and tmr_registers(2)(773)) or                                                       
                            (tmr_registers(0)(773) and tmr_registers(2)(773));                                                         
                                                                                                                                     
        global_tmr_voter(2)(774)  <=    (tmr_registers(0)(774) and tmr_registers(1)(774)) or                                            
                            (tmr_registers(1)(774) and tmr_registers(2)(774)) or                                                       
                            (tmr_registers(0)(774) and tmr_registers(2)(774));                                                         
                                                                                                                                     
        global_tmr_voter(2)(775)  <=    (tmr_registers(0)(775) and tmr_registers(1)(775)) or                                            
                            (tmr_registers(1)(775) and tmr_registers(2)(775)) or                                                       
                            (tmr_registers(0)(775) and tmr_registers(2)(775));                                                         
                                                                                                                                     
        global_tmr_voter(2)(776)  <=    (tmr_registers(0)(776) and tmr_registers(1)(776)) or                                            
                            (tmr_registers(1)(776) and tmr_registers(2)(776)) or                                                       
                            (tmr_registers(0)(776) and tmr_registers(2)(776));                                                         
                                                                                                                                     
        global_tmr_voter(2)(777)  <=    (tmr_registers(0)(777) and tmr_registers(1)(777)) or                                            
                            (tmr_registers(1)(777) and tmr_registers(2)(777)) or                                                       
                            (tmr_registers(0)(777) and tmr_registers(2)(777));                                                         
                                                                                                                                     
        global_tmr_voter(2)(778)  <=    (tmr_registers(0)(778) and tmr_registers(1)(778)) or                                            
                            (tmr_registers(1)(778) and tmr_registers(2)(778)) or                                                       
                            (tmr_registers(0)(778) and tmr_registers(2)(778));                                                         
                                                                                                                                     
        global_tmr_voter(2)(779)  <=    (tmr_registers(0)(779) and tmr_registers(1)(779)) or                                            
                            (tmr_registers(1)(779) and tmr_registers(2)(779)) or                                                       
                            (tmr_registers(0)(779) and tmr_registers(2)(779));                                                         
                                                                                                                                     
        global_tmr_voter(2)(780)  <=    (tmr_registers(0)(780) and tmr_registers(1)(780)) or                                            
                            (tmr_registers(1)(780) and tmr_registers(2)(780)) or                                                       
                            (tmr_registers(0)(780) and tmr_registers(2)(780));                                                         
                                                                                                                                     
        global_tmr_voter(2)(781)  <=    (tmr_registers(0)(781) and tmr_registers(1)(781)) or                                            
                            (tmr_registers(1)(781) and tmr_registers(2)(781)) or                                                       
                            (tmr_registers(0)(781) and tmr_registers(2)(781));                                                         
                                                                                                                                     
        global_tmr_voter(2)(782)  <=    (tmr_registers(0)(782) and tmr_registers(1)(782)) or                                            
                            (tmr_registers(1)(782) and tmr_registers(2)(782)) or                                                       
                            (tmr_registers(0)(782) and tmr_registers(2)(782));                                                         
                                                                                                                                     
        global_tmr_voter(2)(783)  <=    (tmr_registers(0)(783) and tmr_registers(1)(783)) or                                            
                            (tmr_registers(1)(783) and tmr_registers(2)(783)) or                                                       
                            (tmr_registers(0)(783) and tmr_registers(2)(783));                                                         
                                                                                                                                     
        global_tmr_voter(2)(784)  <=    (tmr_registers(0)(784) and tmr_registers(1)(784)) or                                            
                            (tmr_registers(1)(784) and tmr_registers(2)(784)) or                                                       
                            (tmr_registers(0)(784) and tmr_registers(2)(784));                                                         
                                                                                                                                     
        global_tmr_voter(2)(785)  <=    (tmr_registers(0)(785) and tmr_registers(1)(785)) or                                            
                            (tmr_registers(1)(785) and tmr_registers(2)(785)) or                                                       
                            (tmr_registers(0)(785) and tmr_registers(2)(785));                                                         
                                                                                                                                     
        global_tmr_voter(2)(786)  <=    (tmr_registers(0)(786) and tmr_registers(1)(786)) or                                            
                            (tmr_registers(1)(786) and tmr_registers(2)(786)) or                                                       
                            (tmr_registers(0)(786) and tmr_registers(2)(786));                                                         
                                                                                                                                     
        global_tmr_voter(2)(787)  <=    (tmr_registers(0)(787) and tmr_registers(1)(787)) or                                            
                            (tmr_registers(1)(787) and tmr_registers(2)(787)) or                                                       
                            (tmr_registers(0)(787) and tmr_registers(2)(787));                                                         
                                                                                                                                     
        global_tmr_voter(2)(788)  <=    (tmr_registers(0)(788) and tmr_registers(1)(788)) or                                            
                            (tmr_registers(1)(788) and tmr_registers(2)(788)) or                                                       
                            (tmr_registers(0)(788) and tmr_registers(2)(788));                                                         
                                                                                                                                     
        global_tmr_voter(2)(789)  <=    (tmr_registers(0)(789) and tmr_registers(1)(789)) or                                            
                            (tmr_registers(1)(789) and tmr_registers(2)(789)) or                                                       
                            (tmr_registers(0)(789) and tmr_registers(2)(789));                                                         
                                                                                                                                     
        global_tmr_voter(2)(790)  <=    (tmr_registers(0)(790) and tmr_registers(1)(790)) or                                            
                            (tmr_registers(1)(790) and tmr_registers(2)(790)) or                                                       
                            (tmr_registers(0)(790) and tmr_registers(2)(790));                                                         
                                                                                                                                     
        global_tmr_voter(2)(791)  <=    (tmr_registers(0)(791) and tmr_registers(1)(791)) or                                            
                            (tmr_registers(1)(791) and tmr_registers(2)(791)) or                                                       
                            (tmr_registers(0)(791) and tmr_registers(2)(791));                                                         
                                                                                                                                     
        global_tmr_voter(2)(792)  <=    (tmr_registers(0)(792) and tmr_registers(1)(792)) or                                            
                            (tmr_registers(1)(792) and tmr_registers(2)(792)) or                                                       
                            (tmr_registers(0)(792) and tmr_registers(2)(792));                                                         
                                                                                                                                     
        global_tmr_voter(2)(793)  <=    (tmr_registers(0)(793) and tmr_registers(1)(793)) or                                            
                            (tmr_registers(1)(793) and tmr_registers(2)(793)) or                                                       
                            (tmr_registers(0)(793) and tmr_registers(2)(793));                                                         
                                                                                                                                     
        global_tmr_voter(2)(794)  <=    (tmr_registers(0)(794) and tmr_registers(1)(794)) or                                            
                            (tmr_registers(1)(794) and tmr_registers(2)(794)) or                                                       
                            (tmr_registers(0)(794) and tmr_registers(2)(794));                                                         
                                                                                                                                     
        global_tmr_voter(2)(795)  <=    (tmr_registers(0)(795) and tmr_registers(1)(795)) or                                            
                            (tmr_registers(1)(795) and tmr_registers(2)(795)) or                                                       
                            (tmr_registers(0)(795) and tmr_registers(2)(795));                                                         
                                                                                                                                     
        global_tmr_voter(2)(796)  <=    (tmr_registers(0)(796) and tmr_registers(1)(796)) or                                            
                            (tmr_registers(1)(796) and tmr_registers(2)(796)) or                                                       
                            (tmr_registers(0)(796) and tmr_registers(2)(796));                                                         
                                                                                                                                     
        global_tmr_voter(2)(797)  <=    (tmr_registers(0)(797) and tmr_registers(1)(797)) or                                            
                            (tmr_registers(1)(797) and tmr_registers(2)(797)) or                                                       
                            (tmr_registers(0)(797) and tmr_registers(2)(797));                                                         
                                                                                                                                     
        global_tmr_voter(2)(798)  <=    (tmr_registers(0)(798) and tmr_registers(1)(798)) or                                            
                            (tmr_registers(1)(798) and tmr_registers(2)(798)) or                                                       
                            (tmr_registers(0)(798) and tmr_registers(2)(798));                                                         
                                                                                                                                     
        global_tmr_voter(2)(799)  <=    (tmr_registers(0)(799) and tmr_registers(1)(799)) or                                            
                            (tmr_registers(1)(799) and tmr_registers(2)(799)) or                                                       
                            (tmr_registers(0)(799) and tmr_registers(2)(799));                                                         
                                                                                                                                     
        global_tmr_voter(2)(800)  <=    (tmr_registers(0)(800) and tmr_registers(1)(800)) or                                            
                            (tmr_registers(1)(800) and tmr_registers(2)(800)) or                                                       
                            (tmr_registers(0)(800) and tmr_registers(2)(800));                                                         
                                                                                                                                     
        global_tmr_voter(2)(801)  <=    (tmr_registers(0)(801) and tmr_registers(1)(801)) or                                            
                            (tmr_registers(1)(801) and tmr_registers(2)(801)) or                                                       
                            (tmr_registers(0)(801) and tmr_registers(2)(801));                                                         
                                                                                                                                     
        global_tmr_voter(2)(802)  <=    (tmr_registers(0)(802) and tmr_registers(1)(802)) or                                            
                            (tmr_registers(1)(802) and tmr_registers(2)(802)) or                                                       
                            (tmr_registers(0)(802) and tmr_registers(2)(802));                                                         
                                                                                                                                     
        global_tmr_voter(2)(803)  <=    (tmr_registers(0)(803) and tmr_registers(1)(803)) or                                            
                            (tmr_registers(1)(803) and tmr_registers(2)(803)) or                                                       
                            (tmr_registers(0)(803) and tmr_registers(2)(803));                                                         
                                                                                                                                     
        global_tmr_voter(2)(804)  <=    (tmr_registers(0)(804) and tmr_registers(1)(804)) or                                            
                            (tmr_registers(1)(804) and tmr_registers(2)(804)) or                                                       
                            (tmr_registers(0)(804) and tmr_registers(2)(804));                                                         
                                                                                                                                     
        global_tmr_voter(2)(805)  <=    (tmr_registers(0)(805) and tmr_registers(1)(805)) or                                            
                            (tmr_registers(1)(805) and tmr_registers(2)(805)) or                                                       
                            (tmr_registers(0)(805) and tmr_registers(2)(805));                                                         
                                                                                                                                     
        global_tmr_voter(2)(806)  <=    (tmr_registers(0)(806) and tmr_registers(1)(806)) or                                            
                            (tmr_registers(1)(806) and tmr_registers(2)(806)) or                                                       
                            (tmr_registers(0)(806) and tmr_registers(2)(806));                                                         
                                                                                                                                     
        global_tmr_voter(2)(807)  <=    (tmr_registers(0)(807) and tmr_registers(1)(807)) or                                            
                            (tmr_registers(1)(807) and tmr_registers(2)(807)) or                                                       
                            (tmr_registers(0)(807) and tmr_registers(2)(807));                                                         
                                                                                                                                     
        global_tmr_voter(2)(808)  <=    (tmr_registers(0)(808) and tmr_registers(1)(808)) or                                            
                            (tmr_registers(1)(808) and tmr_registers(2)(808)) or                                                       
                            (tmr_registers(0)(808) and tmr_registers(2)(808));                                                         
                                                                                                                                     
        global_tmr_voter(2)(809)  <=    (tmr_registers(0)(809) and tmr_registers(1)(809)) or                                            
                            (tmr_registers(1)(809) and tmr_registers(2)(809)) or                                                       
                            (tmr_registers(0)(809) and tmr_registers(2)(809));                                                         
                                                                                                                                     
        global_tmr_voter(2)(810)  <=    (tmr_registers(0)(810) and tmr_registers(1)(810)) or                                            
                            (tmr_registers(1)(810) and tmr_registers(2)(810)) or                                                       
                            (tmr_registers(0)(810) and tmr_registers(2)(810));                                                         
                                                                                                                                     
        global_tmr_voter(2)(811)  <=    (tmr_registers(0)(811) and tmr_registers(1)(811)) or                                            
                            (tmr_registers(1)(811) and tmr_registers(2)(811)) or                                                       
                            (tmr_registers(0)(811) and tmr_registers(2)(811));                                                         
                                                                                                                                     
        global_tmr_voter(2)(812)  <=    (tmr_registers(0)(812) and tmr_registers(1)(812)) or                                            
                            (tmr_registers(1)(812) and tmr_registers(2)(812)) or                                                       
                            (tmr_registers(0)(812) and tmr_registers(2)(812));                                                         
                                                                                                                                     
        global_tmr_voter(2)(813)  <=    (tmr_registers(0)(813) and tmr_registers(1)(813)) or                                            
                            (tmr_registers(1)(813) and tmr_registers(2)(813)) or                                                       
                            (tmr_registers(0)(813) and tmr_registers(2)(813));                                                         
                                                                                                                                     
        global_tmr_voter(2)(814)  <=    (tmr_registers(0)(814) and tmr_registers(1)(814)) or                                            
                            (tmr_registers(1)(814) and tmr_registers(2)(814)) or                                                       
                            (tmr_registers(0)(814) and tmr_registers(2)(814));                                                         
                                                                                                                                     
        global_tmr_voter(2)(815)  <=    (tmr_registers(0)(815) and tmr_registers(1)(815)) or                                            
                            (tmr_registers(1)(815) and tmr_registers(2)(815)) or                                                       
                            (tmr_registers(0)(815) and tmr_registers(2)(815));                                                         
                                                                                                                                     
        global_tmr_voter(2)(816)  <=    (tmr_registers(0)(816) and tmr_registers(1)(816)) or                                            
                            (tmr_registers(1)(816) and tmr_registers(2)(816)) or                                                       
                            (tmr_registers(0)(816) and tmr_registers(2)(816));                                                         
                                                                                                                                     
        global_tmr_voter(2)(817)  <=    (tmr_registers(0)(817) and tmr_registers(1)(817)) or                                            
                            (tmr_registers(1)(817) and tmr_registers(2)(817)) or                                                       
                            (tmr_registers(0)(817) and tmr_registers(2)(817));                                                         
                                                                                                                                     
        global_tmr_voter(2)(818)  <=    (tmr_registers(0)(818) and tmr_registers(1)(818)) or                                            
                            (tmr_registers(1)(818) and tmr_registers(2)(818)) or                                                       
                            (tmr_registers(0)(818) and tmr_registers(2)(818));                                                         
                                                                                                                                     
        global_tmr_voter(2)(819)  <=    (tmr_registers(0)(819) and tmr_registers(1)(819)) or                                            
                            (tmr_registers(1)(819) and tmr_registers(2)(819)) or                                                       
                            (tmr_registers(0)(819) and tmr_registers(2)(819));                                                         
                                                                                                                                     
        global_tmr_voter(2)(820)  <=    (tmr_registers(0)(820) and tmr_registers(1)(820)) or                                            
                            (tmr_registers(1)(820) and tmr_registers(2)(820)) or                                                       
                            (tmr_registers(0)(820) and tmr_registers(2)(820));                                                         
                                                                                                                                     
        global_tmr_voter(2)(821)  <=    (tmr_registers(0)(821) and tmr_registers(1)(821)) or                                            
                            (tmr_registers(1)(821) and tmr_registers(2)(821)) or                                                       
                            (tmr_registers(0)(821) and tmr_registers(2)(821));                                                         
                                                                                                                                     
        global_tmr_voter(2)(822)  <=    (tmr_registers(0)(822) and tmr_registers(1)(822)) or                                            
                            (tmr_registers(1)(822) and tmr_registers(2)(822)) or                                                       
                            (tmr_registers(0)(822) and tmr_registers(2)(822));                                                         
                                                                                                                                     
        global_tmr_voter(2)(823)  <=    (tmr_registers(0)(823) and tmr_registers(1)(823)) or                                            
                            (tmr_registers(1)(823) and tmr_registers(2)(823)) or                                                       
                            (tmr_registers(0)(823) and tmr_registers(2)(823));                                                         
                                                                                                                                     
        global_tmr_voter(2)(824)  <=    (tmr_registers(0)(824) and tmr_registers(1)(824)) or                                            
                            (tmr_registers(1)(824) and tmr_registers(2)(824)) or                                                       
                            (tmr_registers(0)(824) and tmr_registers(2)(824));                                                         
                                                                                                                                     
        global_tmr_voter(2)(825)  <=    (tmr_registers(0)(825) and tmr_registers(1)(825)) or                                            
                            (tmr_registers(1)(825) and tmr_registers(2)(825)) or                                                       
                            (tmr_registers(0)(825) and tmr_registers(2)(825));                                                         
                                                                                                                                     
        global_tmr_voter(2)(826)  <=    (tmr_registers(0)(826) and tmr_registers(1)(826)) or                                            
                            (tmr_registers(1)(826) and tmr_registers(2)(826)) or                                                       
                            (tmr_registers(0)(826) and tmr_registers(2)(826));                                                         
                                                                                                                                     
        global_tmr_voter(2)(827)  <=    (tmr_registers(0)(827) and tmr_registers(1)(827)) or                                            
                            (tmr_registers(1)(827) and tmr_registers(2)(827)) or                                                       
                            (tmr_registers(0)(827) and tmr_registers(2)(827));                                                         
                                                                                                                                     
        global_tmr_voter(2)(828)  <=    (tmr_registers(0)(828) and tmr_registers(1)(828)) or                                            
                            (tmr_registers(1)(828) and tmr_registers(2)(828)) or                                                       
                            (tmr_registers(0)(828) and tmr_registers(2)(828));                                                         
                                                                                                                                     
        global_tmr_voter(2)(829)  <=    (tmr_registers(0)(829) and tmr_registers(1)(829)) or                                            
                            (tmr_registers(1)(829) and tmr_registers(2)(829)) or                                                       
                            (tmr_registers(0)(829) and tmr_registers(2)(829));                                                         
                                                                                                                                     
        global_tmr_voter(2)(830)  <=    (tmr_registers(0)(830) and tmr_registers(1)(830)) or                                            
                            (tmr_registers(1)(830) and tmr_registers(2)(830)) or                                                       
                            (tmr_registers(0)(830) and tmr_registers(2)(830));                                                         
                                                                                                                                     
        global_tmr_voter(2)(831)  <=    (tmr_registers(0)(831) and tmr_registers(1)(831)) or                                            
                            (tmr_registers(1)(831) and tmr_registers(2)(831)) or                                                       
                            (tmr_registers(0)(831) and tmr_registers(2)(831));                                                         
                                                                                                                                     
        global_tmr_voter(2)(832)  <=    (tmr_registers(0)(832) and tmr_registers(1)(832)) or                                            
                            (tmr_registers(1)(832) and tmr_registers(2)(832)) or                                                       
                            (tmr_registers(0)(832) and tmr_registers(2)(832));                                                         
                                                                                                                                     
        global_tmr_voter(2)(833)  <=    (tmr_registers(0)(833) and tmr_registers(1)(833)) or                                            
                            (tmr_registers(1)(833) and tmr_registers(2)(833)) or                                                       
                            (tmr_registers(0)(833) and tmr_registers(2)(833));                                                         
                                                                                                                                     
        global_tmr_voter(2)(834)  <=    (tmr_registers(0)(834) and tmr_registers(1)(834)) or                                            
                            (tmr_registers(1)(834) and tmr_registers(2)(834)) or                                                       
                            (tmr_registers(0)(834) and tmr_registers(2)(834));                                                         
                                                                                                                                     
        global_tmr_voter(2)(835)  <=    (tmr_registers(0)(835) and tmr_registers(1)(835)) or                                            
                            (tmr_registers(1)(835) and tmr_registers(2)(835)) or                                                       
                            (tmr_registers(0)(835) and tmr_registers(2)(835));                                                         
                                                                                                                                     
        global_tmr_voter(2)(836)  <=    (tmr_registers(0)(836) and tmr_registers(1)(836)) or                                            
                            (tmr_registers(1)(836) and tmr_registers(2)(836)) or                                                       
                            (tmr_registers(0)(836) and tmr_registers(2)(836));                                                         
                                                                                                                                     
        global_tmr_voter(2)(837)  <=    (tmr_registers(0)(837) and tmr_registers(1)(837)) or                                            
                            (tmr_registers(1)(837) and tmr_registers(2)(837)) or                                                       
                            (tmr_registers(0)(837) and tmr_registers(2)(837));                                                         
                                                                                                                                     
        global_tmr_voter(2)(838)  <=    (tmr_registers(0)(838) and tmr_registers(1)(838)) or                                            
                            (tmr_registers(1)(838) and tmr_registers(2)(838)) or                                                       
                            (tmr_registers(0)(838) and tmr_registers(2)(838));                                                         
                                                                                                                                     
        global_tmr_voter(2)(839)  <=    (tmr_registers(0)(839) and tmr_registers(1)(839)) or                                            
                            (tmr_registers(1)(839) and tmr_registers(2)(839)) or                                                       
                            (tmr_registers(0)(839) and tmr_registers(2)(839));                                                         
                                                                                                                                     
        global_tmr_voter(2)(840)  <=    (tmr_registers(0)(840) and tmr_registers(1)(840)) or                                            
                            (tmr_registers(1)(840) and tmr_registers(2)(840)) or                                                       
                            (tmr_registers(0)(840) and tmr_registers(2)(840));                                                         
                                                                                                                                     
        global_tmr_voter(2)(841)  <=    (tmr_registers(0)(841) and tmr_registers(1)(841)) or                                            
                            (tmr_registers(1)(841) and tmr_registers(2)(841)) or                                                       
                            (tmr_registers(0)(841) and tmr_registers(2)(841));                                                         
                                                                                                                                     
        global_tmr_voter(2)(842)  <=    (tmr_registers(0)(842) and tmr_registers(1)(842)) or                                            
                            (tmr_registers(1)(842) and tmr_registers(2)(842)) or                                                       
                            (tmr_registers(0)(842) and tmr_registers(2)(842));                                                         
                                                                                                                                     
        global_tmr_voter(2)(843)  <=    (tmr_registers(0)(843) and tmr_registers(1)(843)) or                                            
                            (tmr_registers(1)(843) and tmr_registers(2)(843)) or                                                       
                            (tmr_registers(0)(843) and tmr_registers(2)(843));                                                         
                                                                                                                                     
        global_tmr_voter(2)(844)  <=    (tmr_registers(0)(844) and tmr_registers(1)(844)) or                                            
                            (tmr_registers(1)(844) and tmr_registers(2)(844)) or                                                       
                            (tmr_registers(0)(844) and tmr_registers(2)(844));                                                         
                                                                                                                                     
        global_tmr_voter(2)(845)  <=    (tmr_registers(0)(845) and tmr_registers(1)(845)) or                                            
                            (tmr_registers(1)(845) and tmr_registers(2)(845)) or                                                       
                            (tmr_registers(0)(845) and tmr_registers(2)(845));                                                         
                                                                                                                                     
        global_tmr_voter(2)(846)  <=    (tmr_registers(0)(846) and tmr_registers(1)(846)) or                                            
                            (tmr_registers(1)(846) and tmr_registers(2)(846)) or                                                       
                            (tmr_registers(0)(846) and tmr_registers(2)(846));                                                         
                                                                                                                                     
        global_tmr_voter(2)(847)  <=    (tmr_registers(0)(847) and tmr_registers(1)(847)) or                                            
                            (tmr_registers(1)(847) and tmr_registers(2)(847)) or                                                       
                            (tmr_registers(0)(847) and tmr_registers(2)(847));                                                         
                                                                                                                                     
        global_tmr_voter(2)(848)  <=    (tmr_registers(0)(848) and tmr_registers(1)(848)) or                                            
                            (tmr_registers(1)(848) and tmr_registers(2)(848)) or                                                       
                            (tmr_registers(0)(848) and tmr_registers(2)(848));                                                         
                                                                                                                                     
        global_tmr_voter(2)(849)  <=    (tmr_registers(0)(849) and tmr_registers(1)(849)) or                                            
                            (tmr_registers(1)(849) and tmr_registers(2)(849)) or                                                       
                            (tmr_registers(0)(849) and tmr_registers(2)(849));                                                         
                                                                                                                                     
        global_tmr_voter(2)(850)  <=    (tmr_registers(0)(850) and tmr_registers(1)(850)) or                                            
                            (tmr_registers(1)(850) and tmr_registers(2)(850)) or                                                       
                            (tmr_registers(0)(850) and tmr_registers(2)(850));                                                         
                                                                                                                                     
        global_tmr_voter(2)(851)  <=    (tmr_registers(0)(851) and tmr_registers(1)(851)) or                                            
                            (tmr_registers(1)(851) and tmr_registers(2)(851)) or                                                       
                            (tmr_registers(0)(851) and tmr_registers(2)(851));                                                         
                                                                                                                                     
        global_tmr_voter(2)(852)  <=    (tmr_registers(0)(852) and tmr_registers(1)(852)) or                                            
                            (tmr_registers(1)(852) and tmr_registers(2)(852)) or                                                       
                            (tmr_registers(0)(852) and tmr_registers(2)(852));                                                         
                                                                                                                                     
        global_tmr_voter(2)(853)  <=    (tmr_registers(0)(853) and tmr_registers(1)(853)) or                                            
                            (tmr_registers(1)(853) and tmr_registers(2)(853)) or                                                       
                            (tmr_registers(0)(853) and tmr_registers(2)(853));                                                         
                                                                                                                                     
        global_tmr_voter(2)(854)  <=    (tmr_registers(0)(854) and tmr_registers(1)(854)) or                                            
                            (tmr_registers(1)(854) and tmr_registers(2)(854)) or                                                       
                            (tmr_registers(0)(854) and tmr_registers(2)(854));                                                         
                                                                                                                                     
        global_tmr_voter(2)(855)  <=    (tmr_registers(0)(855) and tmr_registers(1)(855)) or                                            
                            (tmr_registers(1)(855) and tmr_registers(2)(855)) or                                                       
                            (tmr_registers(0)(855) and tmr_registers(2)(855));                                                         
                                                                                                                                     
        global_tmr_voter(2)(856)  <=    (tmr_registers(0)(856) and tmr_registers(1)(856)) or                                            
                            (tmr_registers(1)(856) and tmr_registers(2)(856)) or                                                       
                            (tmr_registers(0)(856) and tmr_registers(2)(856));                                                         
                                                                                                                                     
        global_tmr_voter(2)(857)  <=    (tmr_registers(0)(857) and tmr_registers(1)(857)) or                                            
                            (tmr_registers(1)(857) and tmr_registers(2)(857)) or                                                       
                            (tmr_registers(0)(857) and tmr_registers(2)(857));                                                         
                                                                                                                                     
        global_tmr_voter(2)(858)  <=    (tmr_registers(0)(858) and tmr_registers(1)(858)) or                                            
                            (tmr_registers(1)(858) and tmr_registers(2)(858)) or                                                       
                            (tmr_registers(0)(858) and tmr_registers(2)(858));                                                         
                                                                                                                                     
        global_tmr_voter(2)(859)  <=    (tmr_registers(0)(859) and tmr_registers(1)(859)) or                                            
                            (tmr_registers(1)(859) and tmr_registers(2)(859)) or                                                       
                            (tmr_registers(0)(859) and tmr_registers(2)(859));                                                         
                                                                                                                                     
        global_tmr_voter(2)(860)  <=    (tmr_registers(0)(860) and tmr_registers(1)(860)) or                                            
                            (tmr_registers(1)(860) and tmr_registers(2)(860)) or                                                       
                            (tmr_registers(0)(860) and tmr_registers(2)(860));                                                         
                                                                                                                                     
        global_tmr_voter(2)(861)  <=    (tmr_registers(0)(861) and tmr_registers(1)(861)) or                                            
                            (tmr_registers(1)(861) and tmr_registers(2)(861)) or                                                       
                            (tmr_registers(0)(861) and tmr_registers(2)(861));                                                         
                                                                                                                                     
        global_tmr_voter(2)(862)  <=    (tmr_registers(0)(862) and tmr_registers(1)(862)) or                                            
                            (tmr_registers(1)(862) and tmr_registers(2)(862)) or                                                       
                            (tmr_registers(0)(862) and tmr_registers(2)(862));                                                         
                                                                                                                                     
        global_tmr_voter(2)(863)  <=    (tmr_registers(0)(863) and tmr_registers(1)(863)) or                                            
                            (tmr_registers(1)(863) and tmr_registers(2)(863)) or                                                       
                            (tmr_registers(0)(863) and tmr_registers(2)(863));                                                         
                                                                                                                                     
        global_tmr_voter(2)(864)  <=    (tmr_registers(0)(864) and tmr_registers(1)(864)) or                                            
                            (tmr_registers(1)(864) and tmr_registers(2)(864)) or                                                       
                            (tmr_registers(0)(864) and tmr_registers(2)(864));                                                         
                                                                                                                                     
        global_tmr_voter(2)(865)  <=    (tmr_registers(0)(865) and tmr_registers(1)(865)) or                                            
                            (tmr_registers(1)(865) and tmr_registers(2)(865)) or                                                       
                            (tmr_registers(0)(865) and tmr_registers(2)(865));                                                         
                                                                                                                                     
        global_tmr_voter(2)(866)  <=    (tmr_registers(0)(866) and tmr_registers(1)(866)) or                                            
                            (tmr_registers(1)(866) and tmr_registers(2)(866)) or                                                       
                            (tmr_registers(0)(866) and tmr_registers(2)(866));                                                         
                                                                                                                                     
        global_tmr_voter(2)(867)  <=    (tmr_registers(0)(867) and tmr_registers(1)(867)) or                                            
                            (tmr_registers(1)(867) and tmr_registers(2)(867)) or                                                       
                            (tmr_registers(0)(867) and tmr_registers(2)(867));                                                         
                                                                                                                                     
        global_tmr_voter(2)(868)  <=    (tmr_registers(0)(868) and tmr_registers(1)(868)) or                                            
                            (tmr_registers(1)(868) and tmr_registers(2)(868)) or                                                       
                            (tmr_registers(0)(868) and tmr_registers(2)(868));                                                         
                                                                                                                                     
        global_tmr_voter(2)(869)  <=    (tmr_registers(0)(869) and tmr_registers(1)(869)) or                                            
                            (tmr_registers(1)(869) and tmr_registers(2)(869)) or                                                       
                            (tmr_registers(0)(869) and tmr_registers(2)(869));                                                         
                                                                                                                                     
        global_tmr_voter(2)(870)  <=    (tmr_registers(0)(870) and tmr_registers(1)(870)) or                                            
                            (tmr_registers(1)(870) and tmr_registers(2)(870)) or                                                       
                            (tmr_registers(0)(870) and tmr_registers(2)(870));                                                         
                                                                                                                                     
        global_tmr_voter(2)(871)  <=    (tmr_registers(0)(871) and tmr_registers(1)(871)) or                                            
                            (tmr_registers(1)(871) and tmr_registers(2)(871)) or                                                       
                            (tmr_registers(0)(871) and tmr_registers(2)(871));                                                         
                                                                                                                                     
        global_tmr_voter(2)(872)  <=    (tmr_registers(0)(872) and tmr_registers(1)(872)) or                                            
                            (tmr_registers(1)(872) and tmr_registers(2)(872)) or                                                       
                            (tmr_registers(0)(872) and tmr_registers(2)(872));                                                         
                                                                                                                                     
        global_tmr_voter(2)(873)  <=    (tmr_registers(0)(873) and tmr_registers(1)(873)) or                                            
                            (tmr_registers(1)(873) and tmr_registers(2)(873)) or                                                       
                            (tmr_registers(0)(873) and tmr_registers(2)(873));                                                         
                                                                                                                                     
        global_tmr_voter(2)(874)  <=    (tmr_registers(0)(874) and tmr_registers(1)(874)) or                                            
                            (tmr_registers(1)(874) and tmr_registers(2)(874)) or                                                       
                            (tmr_registers(0)(874) and tmr_registers(2)(874));                                                         
                                                                                                                                     
        global_tmr_voter(2)(875)  <=    (tmr_registers(0)(875) and tmr_registers(1)(875)) or                                            
                            (tmr_registers(1)(875) and tmr_registers(2)(875)) or                                                       
                            (tmr_registers(0)(875) and tmr_registers(2)(875));                                                         
                                                                                                                                     
        global_tmr_voter(2)(876)  <=    (tmr_registers(0)(876) and tmr_registers(1)(876)) or                                            
                            (tmr_registers(1)(876) and tmr_registers(2)(876)) or                                                       
                            (tmr_registers(0)(876) and tmr_registers(2)(876));                                                         
                                                                                                                                     
        global_tmr_voter(2)(877)  <=    (tmr_registers(0)(877) and tmr_registers(1)(877)) or                                            
                            (tmr_registers(1)(877) and tmr_registers(2)(877)) or                                                       
                            (tmr_registers(0)(877) and tmr_registers(2)(877));                                                         
                                                                                                                                     
        global_tmr_voter(2)(878)  <=    (tmr_registers(0)(878) and tmr_registers(1)(878)) or                                            
                            (tmr_registers(1)(878) and tmr_registers(2)(878)) or                                                       
                            (tmr_registers(0)(878) and tmr_registers(2)(878));                                                         
                                                                                                                                     
        global_tmr_voter(2)(879)  <=    (tmr_registers(0)(879) and tmr_registers(1)(879)) or                                            
                            (tmr_registers(1)(879) and tmr_registers(2)(879)) or                                                       
                            (tmr_registers(0)(879) and tmr_registers(2)(879));                                                         
                                                                                                                                     
        global_tmr_voter(2)(880)  <=    (tmr_registers(0)(880) and tmr_registers(1)(880)) or                                            
                            (tmr_registers(1)(880) and tmr_registers(2)(880)) or                                                       
                            (tmr_registers(0)(880) and tmr_registers(2)(880));                                                         
                                                                                                                                     
        global_tmr_voter(2)(881)  <=    (tmr_registers(0)(881) and tmr_registers(1)(881)) or                                            
                            (tmr_registers(1)(881) and tmr_registers(2)(881)) or                                                       
                            (tmr_registers(0)(881) and tmr_registers(2)(881));                                                         
                                                                                                                                     
        global_tmr_voter(2)(882)  <=    (tmr_registers(0)(882) and tmr_registers(1)(882)) or                                            
                            (tmr_registers(1)(882) and tmr_registers(2)(882)) or                                                       
                            (tmr_registers(0)(882) and tmr_registers(2)(882));                                                         
                                                                                                                                     
        global_tmr_voter(2)(883)  <=    (tmr_registers(0)(883) and tmr_registers(1)(883)) or                                            
                            (tmr_registers(1)(883) and tmr_registers(2)(883)) or                                                       
                            (tmr_registers(0)(883) and tmr_registers(2)(883));                                                         
                                                                                                                                     
        global_tmr_voter(2)(884)  <=    (tmr_registers(0)(884) and tmr_registers(1)(884)) or                                            
                            (tmr_registers(1)(884) and tmr_registers(2)(884)) or                                                       
                            (tmr_registers(0)(884) and tmr_registers(2)(884));                                                         
                                                                                                                                     
        global_tmr_voter(2)(885)  <=    (tmr_registers(0)(885) and tmr_registers(1)(885)) or                                            
                            (tmr_registers(1)(885) and tmr_registers(2)(885)) or                                                       
                            (tmr_registers(0)(885) and tmr_registers(2)(885));                                                         
                                                                                                                                     
        global_tmr_voter(2)(886)  <=    (tmr_registers(0)(886) and tmr_registers(1)(886)) or                                            
                            (tmr_registers(1)(886) and tmr_registers(2)(886)) or                                                       
                            (tmr_registers(0)(886) and tmr_registers(2)(886));                                                         
                                                                                                                                     
        global_tmr_voter(2)(887)  <=    (tmr_registers(0)(887) and tmr_registers(1)(887)) or                                            
                            (tmr_registers(1)(887) and tmr_registers(2)(887)) or                                                       
                            (tmr_registers(0)(887) and tmr_registers(2)(887));                                                         
                                                                                                                                     
        global_tmr_voter(2)(888)  <=    (tmr_registers(0)(888) and tmr_registers(1)(888)) or                                            
                            (tmr_registers(1)(888) and tmr_registers(2)(888)) or                                                       
                            (tmr_registers(0)(888) and tmr_registers(2)(888));                                                         
                                                                                                                                     
        global_tmr_voter(2)(889)  <=    (tmr_registers(0)(889) and tmr_registers(1)(889)) or                                            
                            (tmr_registers(1)(889) and tmr_registers(2)(889)) or                                                       
                            (tmr_registers(0)(889) and tmr_registers(2)(889));                                                         
                                                                                                                                     
        global_tmr_voter(2)(890)  <=    (tmr_registers(0)(890) and tmr_registers(1)(890)) or                                            
                            (tmr_registers(1)(890) and tmr_registers(2)(890)) or                                                       
                            (tmr_registers(0)(890) and tmr_registers(2)(890));                                                         
                                                                                                                                     
        global_tmr_voter(2)(891)  <=    (tmr_registers(0)(891) and tmr_registers(1)(891)) or                                            
                            (tmr_registers(1)(891) and tmr_registers(2)(891)) or                                                       
                            (tmr_registers(0)(891) and tmr_registers(2)(891));                                                         
                                                                                                                                     
        global_tmr_voter(2)(892)  <=    (tmr_registers(0)(892) and tmr_registers(1)(892)) or                                            
                            (tmr_registers(1)(892) and tmr_registers(2)(892)) or                                                       
                            (tmr_registers(0)(892) and tmr_registers(2)(892));                                                         
                                                                                                                                     
        global_tmr_voter(2)(893)  <=    (tmr_registers(0)(893) and tmr_registers(1)(893)) or                                            
                            (tmr_registers(1)(893) and tmr_registers(2)(893)) or                                                       
                            (tmr_registers(0)(893) and tmr_registers(2)(893));                                                         
                                                                                                                                     
        global_tmr_voter(2)(894)  <=    (tmr_registers(0)(894) and tmr_registers(1)(894)) or                                            
                            (tmr_registers(1)(894) and tmr_registers(2)(894)) or                                                       
                            (tmr_registers(0)(894) and tmr_registers(2)(894));                                                         
                                                                                                                                     
        global_tmr_voter(2)(895)  <=    (tmr_registers(0)(895) and tmr_registers(1)(895)) or                                            
                            (tmr_registers(1)(895) and tmr_registers(2)(895)) or                                                       
                            (tmr_registers(0)(895) and tmr_registers(2)(895));                                                         
                                                                                                                                     
        global_tmr_voter(2)(896)  <=    (tmr_registers(0)(896) and tmr_registers(1)(896)) or                                            
                            (tmr_registers(1)(896) and tmr_registers(2)(896)) or                                                       
                            (tmr_registers(0)(896) and tmr_registers(2)(896));                                                         
                                                                                                                                     
        global_tmr_voter(2)(897)  <=    (tmr_registers(0)(897) and tmr_registers(1)(897)) or                                            
                            (tmr_registers(1)(897) and tmr_registers(2)(897)) or                                                       
                            (tmr_registers(0)(897) and tmr_registers(2)(897));                                                         
                                                                                                                                     
        global_tmr_voter(2)(898)  <=    (tmr_registers(0)(898) and tmr_registers(1)(898)) or                                            
                            (tmr_registers(1)(898) and tmr_registers(2)(898)) or                                                       
                            (tmr_registers(0)(898) and tmr_registers(2)(898));                                                         
                                                                                                                                     
        global_tmr_voter(2)(899)  <=    (tmr_registers(0)(899) and tmr_registers(1)(899)) or                                            
                            (tmr_registers(1)(899) and tmr_registers(2)(899)) or                                                       
                            (tmr_registers(0)(899) and tmr_registers(2)(899));                                                         
                                                                                                                                     
        global_tmr_voter(2)(900)  <=    (tmr_registers(0)(900) and tmr_registers(1)(900)) or                                            
                            (tmr_registers(1)(900) and tmr_registers(2)(900)) or                                                       
                            (tmr_registers(0)(900) and tmr_registers(2)(900));                                                         
                                                                                                                                     
        global_tmr_voter(2)(901)  <=    (tmr_registers(0)(901) and tmr_registers(1)(901)) or                                            
                            (tmr_registers(1)(901) and tmr_registers(2)(901)) or                                                       
                            (tmr_registers(0)(901) and tmr_registers(2)(901));                                                         
                                                                                                                                     
        global_tmr_voter(2)(902)  <=    (tmr_registers(0)(902) and tmr_registers(1)(902)) or                                            
                            (tmr_registers(1)(902) and tmr_registers(2)(902)) or                                                       
                            (tmr_registers(0)(902) and tmr_registers(2)(902));                                                         
                                                                                                                                     
        global_tmr_voter(2)(903)  <=    (tmr_registers(0)(903) and tmr_registers(1)(903)) or                                            
                            (tmr_registers(1)(903) and tmr_registers(2)(903)) or                                                       
                            (tmr_registers(0)(903) and tmr_registers(2)(903));                                                         
                                                                                                                                     
        global_tmr_voter(2)(904)  <=    (tmr_registers(0)(904) and tmr_registers(1)(904)) or                                            
                            (tmr_registers(1)(904) and tmr_registers(2)(904)) or                                                       
                            (tmr_registers(0)(904) and tmr_registers(2)(904));                                                         
                                                                                                                                     
        global_tmr_voter(2)(905)  <=    (tmr_registers(0)(905) and tmr_registers(1)(905)) or                                            
                            (tmr_registers(1)(905) and tmr_registers(2)(905)) or                                                       
                            (tmr_registers(0)(905) and tmr_registers(2)(905));                                                         
                                                                                                                                     
        global_tmr_voter(2)(906)  <=    (tmr_registers(0)(906) and tmr_registers(1)(906)) or                                            
                            (tmr_registers(1)(906) and tmr_registers(2)(906)) or                                                       
                            (tmr_registers(0)(906) and tmr_registers(2)(906));                                                         
                                                                                                                                     
        global_tmr_voter(2)(907)  <=    (tmr_registers(0)(907) and tmr_registers(1)(907)) or                                            
                            (tmr_registers(1)(907) and tmr_registers(2)(907)) or                                                       
                            (tmr_registers(0)(907) and tmr_registers(2)(907));                                                         
                                                                                                                                     
        global_tmr_voter(2)(908)  <=    (tmr_registers(0)(908) and tmr_registers(1)(908)) or                                            
                            (tmr_registers(1)(908) and tmr_registers(2)(908)) or                                                       
                            (tmr_registers(0)(908) and tmr_registers(2)(908));                                                         
                                                                                                                                     
        global_tmr_voter(2)(909)  <=    (tmr_registers(0)(909) and tmr_registers(1)(909)) or                                            
                            (tmr_registers(1)(909) and tmr_registers(2)(909)) or                                                       
                            (tmr_registers(0)(909) and tmr_registers(2)(909));                                                         
                                                                                                                                     
        global_tmr_voter(2)(910)  <=    (tmr_registers(0)(910) and tmr_registers(1)(910)) or                                            
                            (tmr_registers(1)(910) and tmr_registers(2)(910)) or                                                       
                            (tmr_registers(0)(910) and tmr_registers(2)(910));                                                         
                                                                                                                                     
        global_tmr_voter(2)(911)  <=    (tmr_registers(0)(911) and tmr_registers(1)(911)) or                                            
                            (tmr_registers(1)(911) and tmr_registers(2)(911)) or                                                       
                            (tmr_registers(0)(911) and tmr_registers(2)(911));                                                         
                                                                                                                                     
        global_tmr_voter(2)(912)  <=    (tmr_registers(0)(912) and tmr_registers(1)(912)) or                                            
                            (tmr_registers(1)(912) and tmr_registers(2)(912)) or                                                       
                            (tmr_registers(0)(912) and tmr_registers(2)(912));                                                         
                                                                                                                                     
        global_tmr_voter(2)(913)  <=    (tmr_registers(0)(913) and tmr_registers(1)(913)) or                                            
                            (tmr_registers(1)(913) and tmr_registers(2)(913)) or                                                       
                            (tmr_registers(0)(913) and tmr_registers(2)(913));                                                         
                                                                                                                                     
        global_tmr_voter(2)(914)  <=    (tmr_registers(0)(914) and tmr_registers(1)(914)) or                                            
                            (tmr_registers(1)(914) and tmr_registers(2)(914)) or                                                       
                            (tmr_registers(0)(914) and tmr_registers(2)(914));                                                         
                                                                                                                                     
        global_tmr_voter(2)(915)  <=    (tmr_registers(0)(915) and tmr_registers(1)(915)) or                                            
                            (tmr_registers(1)(915) and tmr_registers(2)(915)) or                                                       
                            (tmr_registers(0)(915) and tmr_registers(2)(915));                                                         
                                                                                                                                     
        global_tmr_voter(2)(916)  <=    (tmr_registers(0)(916) and tmr_registers(1)(916)) or                                            
                            (tmr_registers(1)(916) and tmr_registers(2)(916)) or                                                       
                            (tmr_registers(0)(916) and tmr_registers(2)(916));                                                         
                                                                                                                                     
        global_tmr_voter(2)(917)  <=    (tmr_registers(0)(917) and tmr_registers(1)(917)) or                                            
                            (tmr_registers(1)(917) and tmr_registers(2)(917)) or                                                       
                            (tmr_registers(0)(917) and tmr_registers(2)(917));                                                         
                                                                                                                                     
        global_tmr_voter(2)(918)  <=    (tmr_registers(0)(918) and tmr_registers(1)(918)) or                                            
                            (tmr_registers(1)(918) and tmr_registers(2)(918)) or                                                       
                            (tmr_registers(0)(918) and tmr_registers(2)(918));                                                         
                                                                                                                                     
        global_tmr_voter(2)(919)  <=    (tmr_registers(0)(919) and tmr_registers(1)(919)) or                                            
                            (tmr_registers(1)(919) and tmr_registers(2)(919)) or                                                       
                            (tmr_registers(0)(919) and tmr_registers(2)(919));                                                         
                                                                                                                                     
        global_tmr_voter(2)(920)  <=    (tmr_registers(0)(920) and tmr_registers(1)(920)) or                                            
                            (tmr_registers(1)(920) and tmr_registers(2)(920)) or                                                       
                            (tmr_registers(0)(920) and tmr_registers(2)(920));                                                         
                                                                                                                                     
        global_tmr_voter(2)(921)  <=    (tmr_registers(0)(921) and tmr_registers(1)(921)) or                                            
                            (tmr_registers(1)(921) and tmr_registers(2)(921)) or                                                       
                            (tmr_registers(0)(921) and tmr_registers(2)(921));                                                         
                                                                                                                                     
        global_tmr_voter(2)(922)  <=    (tmr_registers(0)(922) and tmr_registers(1)(922)) or                                            
                            (tmr_registers(1)(922) and tmr_registers(2)(922)) or                                                       
                            (tmr_registers(0)(922) and tmr_registers(2)(922));                                                         
                                                                                                                                     
        global_tmr_voter(2)(923)  <=    (tmr_registers(0)(923) and tmr_registers(1)(923)) or                                            
                            (tmr_registers(1)(923) and tmr_registers(2)(923)) or                                                       
                            (tmr_registers(0)(923) and tmr_registers(2)(923));                                                         
                                                                                                                                     
        global_tmr_voter(2)(924)  <=    (tmr_registers(0)(924) and tmr_registers(1)(924)) or                                            
                            (tmr_registers(1)(924) and tmr_registers(2)(924)) or                                                       
                            (tmr_registers(0)(924) and tmr_registers(2)(924));                                                         
                                                                                                                                     
        global_tmr_voter(2)(925)  <=    (tmr_registers(0)(925) and tmr_registers(1)(925)) or                                            
                            (tmr_registers(1)(925) and tmr_registers(2)(925)) or                                                       
                            (tmr_registers(0)(925) and tmr_registers(2)(925));                                                         
                                                                                                                                     
        global_tmr_voter(2)(926)  <=    (tmr_registers(0)(926) and tmr_registers(1)(926)) or                                            
                            (tmr_registers(1)(926) and tmr_registers(2)(926)) or                                                       
                            (tmr_registers(0)(926) and tmr_registers(2)(926));                                                         
                                                                                                                                     
        global_tmr_voter(2)(927)  <=    (tmr_registers(0)(927) and tmr_registers(1)(927)) or                                            
                            (tmr_registers(1)(927) and tmr_registers(2)(927)) or                                                       
                            (tmr_registers(0)(927) and tmr_registers(2)(927));                                                         
                                                                                                                                     
        global_tmr_voter(2)(928)  <=    (tmr_registers(0)(928) and tmr_registers(1)(928)) or                                            
                            (tmr_registers(1)(928) and tmr_registers(2)(928)) or                                                       
                            (tmr_registers(0)(928) and tmr_registers(2)(928));                                                         
                                                                                                                                     
        global_tmr_voter(2)(929)  <=    (tmr_registers(0)(929) and tmr_registers(1)(929)) or                                            
                            (tmr_registers(1)(929) and tmr_registers(2)(929)) or                                                       
                            (tmr_registers(0)(929) and tmr_registers(2)(929));                                                         
                                                                                                                                     
        global_tmr_voter(2)(930)  <=    (tmr_registers(0)(930) and tmr_registers(1)(930)) or                                            
                            (tmr_registers(1)(930) and tmr_registers(2)(930)) or                                                       
                            (tmr_registers(0)(930) and tmr_registers(2)(930));                                                         
                                                                                                                                     
        global_tmr_voter(2)(931)  <=    (tmr_registers(0)(931) and tmr_registers(1)(931)) or                                            
                            (tmr_registers(1)(931) and tmr_registers(2)(931)) or                                                       
                            (tmr_registers(0)(931) and tmr_registers(2)(931));                                                         
                                                                                                                                     
        global_tmr_voter(2)(932)  <=    (tmr_registers(0)(932) and tmr_registers(1)(932)) or                                            
                            (tmr_registers(1)(932) and tmr_registers(2)(932)) or                                                       
                            (tmr_registers(0)(932) and tmr_registers(2)(932));                                                         
                                                                                                                                     
        global_tmr_voter(2)(933)  <=    (tmr_registers(0)(933) and tmr_registers(1)(933)) or                                            
                            (tmr_registers(1)(933) and tmr_registers(2)(933)) or                                                       
                            (tmr_registers(0)(933) and tmr_registers(2)(933));                                                         
                                                                                                                                     
        global_tmr_voter(2)(934)  <=    (tmr_registers(0)(934) and tmr_registers(1)(934)) or                                            
                            (tmr_registers(1)(934) and tmr_registers(2)(934)) or                                                       
                            (tmr_registers(0)(934) and tmr_registers(2)(934));                                                         
                                                                                                                                     
        global_tmr_voter(2)(935)  <=    (tmr_registers(0)(935) and tmr_registers(1)(935)) or                                            
                            (tmr_registers(1)(935) and tmr_registers(2)(935)) or                                                       
                            (tmr_registers(0)(935) and tmr_registers(2)(935));                                                         
                                                                                                                                     
        global_tmr_voter(2)(936)  <=    (tmr_registers(0)(936) and tmr_registers(1)(936)) or                                            
                            (tmr_registers(1)(936) and tmr_registers(2)(936)) or                                                       
                            (tmr_registers(0)(936) and tmr_registers(2)(936));                                                         
                                                                                                                                     
        global_tmr_voter(2)(937)  <=    (tmr_registers(0)(937) and tmr_registers(1)(937)) or                                            
                            (tmr_registers(1)(937) and tmr_registers(2)(937)) or                                                       
                            (tmr_registers(0)(937) and tmr_registers(2)(937));                                                         
                                                                                                                                     
        global_tmr_voter(2)(938)  <=    (tmr_registers(0)(938) and tmr_registers(1)(938)) or                                            
                            (tmr_registers(1)(938) and tmr_registers(2)(938)) or                                                       
                            (tmr_registers(0)(938) and tmr_registers(2)(938));                                                         
                                                                                                                                     
        global_tmr_voter(2)(939)  <=    (tmr_registers(0)(939) and tmr_registers(1)(939)) or                                            
                            (tmr_registers(1)(939) and tmr_registers(2)(939)) or                                                       
                            (tmr_registers(0)(939) and tmr_registers(2)(939));                                                         
                                                                                                                                     
        global_tmr_voter(2)(940)  <=    (tmr_registers(0)(940) and tmr_registers(1)(940)) or                                            
                            (tmr_registers(1)(940) and tmr_registers(2)(940)) or                                                       
                            (tmr_registers(0)(940) and tmr_registers(2)(940));                                                         
                                                                                                                                     
        global_tmr_voter(2)(941)  <=    (tmr_registers(0)(941) and tmr_registers(1)(941)) or                                            
                            (tmr_registers(1)(941) and tmr_registers(2)(941)) or                                                       
                            (tmr_registers(0)(941) and tmr_registers(2)(941));                                                         
                                                                                                                                     
        global_tmr_voter(2)(942)  <=    (tmr_registers(0)(942) and tmr_registers(1)(942)) or                                            
                            (tmr_registers(1)(942) and tmr_registers(2)(942)) or                                                       
                            (tmr_registers(0)(942) and tmr_registers(2)(942));                                                         
                                                                                                                                     
        global_tmr_voter(2)(943)  <=    (tmr_registers(0)(943) and tmr_registers(1)(943)) or                                            
                            (tmr_registers(1)(943) and tmr_registers(2)(943)) or                                                       
                            (tmr_registers(0)(943) and tmr_registers(2)(943));                                                         
                                                                                                                                     
        global_tmr_voter(2)(944)  <=    (tmr_registers(0)(944) and tmr_registers(1)(944)) or                                            
                            (tmr_registers(1)(944) and tmr_registers(2)(944)) or                                                       
                            (tmr_registers(0)(944) and tmr_registers(2)(944));                                                         
                                                                                                                                     
        global_tmr_voter(2)(945)  <=    (tmr_registers(0)(945) and tmr_registers(1)(945)) or                                            
                            (tmr_registers(1)(945) and tmr_registers(2)(945)) or                                                       
                            (tmr_registers(0)(945) and tmr_registers(2)(945));                                                         
                                                                                                                                     
        global_tmr_voter(2)(946)  <=    (tmr_registers(0)(946) and tmr_registers(1)(946)) or                                            
                            (tmr_registers(1)(946) and tmr_registers(2)(946)) or                                                       
                            (tmr_registers(0)(946) and tmr_registers(2)(946));                                                         
                                                                                                                                     
        global_tmr_voter(2)(947)  <=    (tmr_registers(0)(947) and tmr_registers(1)(947)) or                                            
                            (tmr_registers(1)(947) and tmr_registers(2)(947)) or                                                       
                            (tmr_registers(0)(947) and tmr_registers(2)(947));                                                         
                                                                                                                                     
        global_tmr_voter(2)(948)  <=    (tmr_registers(0)(948) and tmr_registers(1)(948)) or                                            
                            (tmr_registers(1)(948) and tmr_registers(2)(948)) or                                                       
                            (tmr_registers(0)(948) and tmr_registers(2)(948));                                                         
                                                                                                                                     
        global_tmr_voter(2)(949)  <=    (tmr_registers(0)(949) and tmr_registers(1)(949)) or                                            
                            (tmr_registers(1)(949) and tmr_registers(2)(949)) or                                                       
                            (tmr_registers(0)(949) and tmr_registers(2)(949));                                                         
                                                                                                                                     
        global_tmr_voter(2)(950)  <=    (tmr_registers(0)(950) and tmr_registers(1)(950)) or                                            
                            (tmr_registers(1)(950) and tmr_registers(2)(950)) or                                                       
                            (tmr_registers(0)(950) and tmr_registers(2)(950));                                                         
                                                                                                                                     
        global_tmr_voter(2)(951)  <=    (tmr_registers(0)(951) and tmr_registers(1)(951)) or                                            
                            (tmr_registers(1)(951) and tmr_registers(2)(951)) or                                                       
                            (tmr_registers(0)(951) and tmr_registers(2)(951));                                                         
                                                                                                                                     
        global_tmr_voter(2)(952)  <=    (tmr_registers(0)(952) and tmr_registers(1)(952)) or                                            
                            (tmr_registers(1)(952) and tmr_registers(2)(952)) or                                                       
                            (tmr_registers(0)(952) and tmr_registers(2)(952));                                                         
                                                                                                                                     
        global_tmr_voter(2)(953)  <=    (tmr_registers(0)(953) and tmr_registers(1)(953)) or                                            
                            (tmr_registers(1)(953) and tmr_registers(2)(953)) or                                                       
                            (tmr_registers(0)(953) and tmr_registers(2)(953));                                                         
                                                                                                                                     
        global_tmr_voter(2)(954)  <=    (tmr_registers(0)(954) and tmr_registers(1)(954)) or                                            
                            (tmr_registers(1)(954) and tmr_registers(2)(954)) or                                                       
                            (tmr_registers(0)(954) and tmr_registers(2)(954));                                                         
                                                                                                                                     
        global_tmr_voter(2)(955)  <=    (tmr_registers(0)(955) and tmr_registers(1)(955)) or                                            
                            (tmr_registers(1)(955) and tmr_registers(2)(955)) or                                                       
                            (tmr_registers(0)(955) and tmr_registers(2)(955));                                                         
                                                                                                                                     
        global_tmr_voter(2)(956)  <=    (tmr_registers(0)(956) and tmr_registers(1)(956)) or                                            
                            (tmr_registers(1)(956) and tmr_registers(2)(956)) or                                                       
                            (tmr_registers(0)(956) and tmr_registers(2)(956));                                                         
                                                                                                                                     
        global_tmr_voter(2)(957)  <=    (tmr_registers(0)(957) and tmr_registers(1)(957)) or                                            
                            (tmr_registers(1)(957) and tmr_registers(2)(957)) or                                                       
                            (tmr_registers(0)(957) and tmr_registers(2)(957));                                                         
                                                                                                                                     
        global_tmr_voter(2)(958)  <=    (tmr_registers(0)(958) and tmr_registers(1)(958)) or                                            
                            (tmr_registers(1)(958) and tmr_registers(2)(958)) or                                                       
                            (tmr_registers(0)(958) and tmr_registers(2)(958));                                                         
                                                                                                                                     
        global_tmr_voter(2)(959)  <=    (tmr_registers(0)(959) and tmr_registers(1)(959)) or                                            
                            (tmr_registers(1)(959) and tmr_registers(2)(959)) or                                                       
                            (tmr_registers(0)(959) and tmr_registers(2)(959));                                                         
                                                                                                                                     
        global_tmr_voter(2)(960)  <=    (tmr_registers(0)(960) and tmr_registers(1)(960)) or                                            
                            (tmr_registers(1)(960) and tmr_registers(2)(960)) or                                                       
                            (tmr_registers(0)(960) and tmr_registers(2)(960));                                                         
                                                                                                                                     
        global_tmr_voter(2)(961)  <=    (tmr_registers(0)(961) and tmr_registers(1)(961)) or                                            
                            (tmr_registers(1)(961) and tmr_registers(2)(961)) or                                                       
                            (tmr_registers(0)(961) and tmr_registers(2)(961));                                                         
                                                                                                                                     
        global_tmr_voter(2)(962)  <=    (tmr_registers(0)(962) and tmr_registers(1)(962)) or                                            
                            (tmr_registers(1)(962) and tmr_registers(2)(962)) or                                                       
                            (tmr_registers(0)(962) and tmr_registers(2)(962));                                                         
                                                                                                                                     
        global_tmr_voter(2)(963)  <=    (tmr_registers(0)(963) and tmr_registers(1)(963)) or                                            
                            (tmr_registers(1)(963) and tmr_registers(2)(963)) or                                                       
                            (tmr_registers(0)(963) and tmr_registers(2)(963));                                                         
                                                                                                                                     
        global_tmr_voter(2)(964)  <=    (tmr_registers(0)(964) and tmr_registers(1)(964)) or                                            
                            (tmr_registers(1)(964) and tmr_registers(2)(964)) or                                                       
                            (tmr_registers(0)(964) and tmr_registers(2)(964));                                                         
                                                                                                                                     
        global_tmr_voter(2)(965)  <=    (tmr_registers(0)(965) and tmr_registers(1)(965)) or                                            
                            (tmr_registers(1)(965) and tmr_registers(2)(965)) or                                                       
                            (tmr_registers(0)(965) and tmr_registers(2)(965));                                                         
                                                                                                                                     
        global_tmr_voter(2)(966)  <=    (tmr_registers(0)(966) and tmr_registers(1)(966)) or                                            
                            (tmr_registers(1)(966) and tmr_registers(2)(966)) or                                                       
                            (tmr_registers(0)(966) and tmr_registers(2)(966));                                                         
                                                                                                                                     
        global_tmr_voter(2)(967)  <=    (tmr_registers(0)(967) and tmr_registers(1)(967)) or                                            
                            (tmr_registers(1)(967) and tmr_registers(2)(967)) or                                                       
                            (tmr_registers(0)(967) and tmr_registers(2)(967));                                                         
                                                                                                                                     
        global_tmr_voter(2)(968)  <=    (tmr_registers(0)(968) and tmr_registers(1)(968)) or                                            
                            (tmr_registers(1)(968) and tmr_registers(2)(968)) or                                                       
                            (tmr_registers(0)(968) and tmr_registers(2)(968));                                                         
                                                                                                                                     
        global_tmr_voter(2)(969)  <=    (tmr_registers(0)(969) and tmr_registers(1)(969)) or                                            
                            (tmr_registers(1)(969) and tmr_registers(2)(969)) or                                                       
                            (tmr_registers(0)(969) and tmr_registers(2)(969));                                                         
                                                                                                                                     
        global_tmr_voter(2)(970)  <=    (tmr_registers(0)(970) and tmr_registers(1)(970)) or                                            
                            (tmr_registers(1)(970) and tmr_registers(2)(970)) or                                                       
                            (tmr_registers(0)(970) and tmr_registers(2)(970));                                                         
                                                                                                                                     
        global_tmr_voter(2)(971)  <=    (tmr_registers(0)(971) and tmr_registers(1)(971)) or                                            
                            (tmr_registers(1)(971) and tmr_registers(2)(971)) or                                                       
                            (tmr_registers(0)(971) and tmr_registers(2)(971));                                                         
                                                                                                                                     
        global_tmr_voter(2)(972)  <=    (tmr_registers(0)(972) and tmr_registers(1)(972)) or                                            
                            (tmr_registers(1)(972) and tmr_registers(2)(972)) or                                                       
                            (tmr_registers(0)(972) and tmr_registers(2)(972));                                                         
                                                                                                                                     
        global_tmr_voter(2)(973)  <=    (tmr_registers(0)(973) and tmr_registers(1)(973)) or                                            
                            (tmr_registers(1)(973) and tmr_registers(2)(973)) or                                                       
                            (tmr_registers(0)(973) and tmr_registers(2)(973));                                                         
                                                                                                                                     
        global_tmr_voter(2)(974)  <=    (tmr_registers(0)(974) and tmr_registers(1)(974)) or                                            
                            (tmr_registers(1)(974) and tmr_registers(2)(974)) or                                                       
                            (tmr_registers(0)(974) and tmr_registers(2)(974));                                                         
                                                                                                                                     
        global_tmr_voter(2)(975)  <=    (tmr_registers(0)(975) and tmr_registers(1)(975)) or                                            
                            (tmr_registers(1)(975) and tmr_registers(2)(975)) or                                                       
                            (tmr_registers(0)(975) and tmr_registers(2)(975));                                                         
                                                                                                                                     
        global_tmr_voter(2)(976)  <=    (tmr_registers(0)(976) and tmr_registers(1)(976)) or                                            
                            (tmr_registers(1)(976) and tmr_registers(2)(976)) or                                                       
                            (tmr_registers(0)(976) and tmr_registers(2)(976));                                                         
                                                                                                                                     
        global_tmr_voter(2)(977)  <=    (tmr_registers(0)(977) and tmr_registers(1)(977)) or                                            
                            (tmr_registers(1)(977) and tmr_registers(2)(977)) or                                                       
                            (tmr_registers(0)(977) and tmr_registers(2)(977));                                                         
                                                                                                                                     
        global_tmr_voter(2)(978)  <=    (tmr_registers(0)(978) and tmr_registers(1)(978)) or                                            
                            (tmr_registers(1)(978) and tmr_registers(2)(978)) or                                                       
                            (tmr_registers(0)(978) and tmr_registers(2)(978));                                                         
                                                                                                                                     
        global_tmr_voter(2)(979)  <=    (tmr_registers(0)(979) and tmr_registers(1)(979)) or                                            
                            (tmr_registers(1)(979) and tmr_registers(2)(979)) or                                                       
                            (tmr_registers(0)(979) and tmr_registers(2)(979));                                                         
                                                                                                                                     
        global_tmr_voter(2)(980)  <=    (tmr_registers(0)(980) and tmr_registers(1)(980)) or                                            
                            (tmr_registers(1)(980) and tmr_registers(2)(980)) or                                                       
                            (tmr_registers(0)(980) and tmr_registers(2)(980));                                                         
                                                                                                                                     
        global_tmr_voter(2)(981)  <=    (tmr_registers(0)(981) and tmr_registers(1)(981)) or                                            
                            (tmr_registers(1)(981) and tmr_registers(2)(981)) or                                                       
                            (tmr_registers(0)(981) and tmr_registers(2)(981));                                                         
                                                                                                                                     
        global_tmr_voter(2)(982)  <=    (tmr_registers(0)(982) and tmr_registers(1)(982)) or                                            
                            (tmr_registers(1)(982) and tmr_registers(2)(982)) or                                                       
                            (tmr_registers(0)(982) and tmr_registers(2)(982));                                                         
                                                                                                                                     
        global_tmr_voter(2)(983)  <=    (tmr_registers(0)(983) and tmr_registers(1)(983)) or                                            
                            (tmr_registers(1)(983) and tmr_registers(2)(983)) or                                                       
                            (tmr_registers(0)(983) and tmr_registers(2)(983));                                                         
                                                                                                                                     
        global_tmr_voter(2)(984)  <=    (tmr_registers(0)(984) and tmr_registers(1)(984)) or                                            
                            (tmr_registers(1)(984) and tmr_registers(2)(984)) or                                                       
                            (tmr_registers(0)(984) and tmr_registers(2)(984));                                                         
                                                                                                                                     
        global_tmr_voter(2)(985)  <=    (tmr_registers(0)(985) and tmr_registers(1)(985)) or                                            
                            (tmr_registers(1)(985) and tmr_registers(2)(985)) or                                                       
                            (tmr_registers(0)(985) and tmr_registers(2)(985));                                                         
                                                                                                                                     
        global_tmr_voter(2)(986)  <=    (tmr_registers(0)(986) and tmr_registers(1)(986)) or                                            
                            (tmr_registers(1)(986) and tmr_registers(2)(986)) or                                                       
                            (tmr_registers(0)(986) and tmr_registers(2)(986));                                                         
                                                                                                                                     
        global_tmr_voter(2)(987)  <=    (tmr_registers(0)(987) and tmr_registers(1)(987)) or                                            
                            (tmr_registers(1)(987) and tmr_registers(2)(987)) or                                                       
                            (tmr_registers(0)(987) and tmr_registers(2)(987));                                                         
                                                                                                                                     
        global_tmr_voter(2)(988)  <=    (tmr_registers(0)(988) and tmr_registers(1)(988)) or                                            
                            (tmr_registers(1)(988) and tmr_registers(2)(988)) or                                                       
                            (tmr_registers(0)(988) and tmr_registers(2)(988));                                                         
                                                                                                                                     
        global_tmr_voter(2)(989)  <=    (tmr_registers(0)(989) and tmr_registers(1)(989)) or                                            
                            (tmr_registers(1)(989) and tmr_registers(2)(989)) or                                                       
                            (tmr_registers(0)(989) and tmr_registers(2)(989));                                                         
                                                                                                                                     
        global_tmr_voter(2)(990)  <=    (tmr_registers(0)(990) and tmr_registers(1)(990)) or                                            
                            (tmr_registers(1)(990) and tmr_registers(2)(990)) or                                                       
                            (tmr_registers(0)(990) and tmr_registers(2)(990));                                                         
                                                                                                                                     
        global_tmr_voter(2)(991)  <=    (tmr_registers(0)(991) and tmr_registers(1)(991)) or                                            
                            (tmr_registers(1)(991) and tmr_registers(2)(991)) or                                                       
                            (tmr_registers(0)(991) and tmr_registers(2)(991));                                                         
                                                                                                                                     
        global_tmr_voter(2)(992)  <=    (tmr_registers(0)(992) and tmr_registers(1)(992)) or                                            
                            (tmr_registers(1)(992) and tmr_registers(2)(992)) or                                                       
                            (tmr_registers(0)(992) and tmr_registers(2)(992));                                                         
                                                                                                                                     
        global_tmr_voter(2)(993)  <=    (tmr_registers(0)(993) and tmr_registers(1)(993)) or                                            
                            (tmr_registers(1)(993) and tmr_registers(2)(993)) or                                                       
                            (tmr_registers(0)(993) and tmr_registers(2)(993));                                                         
                                                                                                                                     
        global_tmr_voter(2)(994)  <=    (tmr_registers(0)(994) and tmr_registers(1)(994)) or                                            
                            (tmr_registers(1)(994) and tmr_registers(2)(994)) or                                                       
                            (tmr_registers(0)(994) and tmr_registers(2)(994));                                                         
                                                                                                                                     
        global_tmr_voter(2)(995)  <=    (tmr_registers(0)(995) and tmr_registers(1)(995)) or                                            
                            (tmr_registers(1)(995) and tmr_registers(2)(995)) or                                                       
                            (tmr_registers(0)(995) and tmr_registers(2)(995));                                                         
                                                                                                                                     
        global_tmr_voter(2)(996)  <=    (tmr_registers(0)(996) and tmr_registers(1)(996)) or                                            
                            (tmr_registers(1)(996) and tmr_registers(2)(996)) or                                                       
                            (tmr_registers(0)(996) and tmr_registers(2)(996));                                                         
                                                                                                                                     
        global_tmr_voter(2)(997)  <=    (tmr_registers(0)(997) and tmr_registers(1)(997)) or                                            
                            (tmr_registers(1)(997) and tmr_registers(2)(997)) or                                                       
                            (tmr_registers(0)(997) and tmr_registers(2)(997));                                                         
                                                                                                                                     
        global_tmr_voter(2)(998)  <=    (tmr_registers(0)(998) and tmr_registers(1)(998)) or                                            
                            (tmr_registers(1)(998) and tmr_registers(2)(998)) or                                                       
                            (tmr_registers(0)(998) and tmr_registers(2)(998));                                                         
                                                                                                                                     
        global_tmr_voter(2)(999)  <=    (tmr_registers(0)(999) and tmr_registers(1)(999)) or                                            
                            (tmr_registers(1)(999) and tmr_registers(2)(999)) or                                                       
                            (tmr_registers(0)(999) and tmr_registers(2)(999));                                                         
                                                                                                                                         
    ------------------------------------------                                                                                           
    -- Outputs                                                                                                                           
    ------------------------------------------                                                                                           
                                                                                                                                         
    data_out(0) <= global_tmr_voter(0)(nb_reg-4);                                                                                        
    data_out(1) <= global_tmr_voter(1)(nb_reg-3);                                                                                        
    data_out(2) <= global_tmr_voter(2)(nb_reg-2);                                                                                        
    data_out(3) <= '0';                                                                                                                
                                                                                                                                         
                                                                                                                                         
end generate GLOBAL_TMR_MITIGATION;                                                                                                      
                                                                                                                                         
                                                                                                                                         
end rtl;                                                                                                                                 
