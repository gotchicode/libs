library IEEE;                                                                                            
use IEEE.std_logic_1164.all;                                                                             
use IEEE.numeric_std.all;                                                                                
use     ieee.math_real.all;                                                                              
                                                                                                         
entity fir_with_tree is                                                                                            
 port (                                                                                                  
            clk             : in std_logic;                                                              
                                                                                                         
            data_in         : in std_logic_vector(11 downto 0);                                          
            data_in_en      : in std_logic;                                                              
                                                                                                         
			data_out		: out std_logic_vector(11 downto 0);                                          
			data_out_en		: out std_logic                                                               
                                                                                                         
 );                                                                                                      
end entity fir_with_tree;                                                                                          
                                                                                                         
architecture rtl of fir_with_tree is                                                                               
                                                                                                         
                                                                                                         
                                                                                                         
constant nb_taps                        : integer:=2048;                                                   
type taps_type                          is array (0 to nb_taps-1) of signed(13 downto 0);                
signal taps                             : taps_type;                                                     
type fir_reg_type                       is array (0 to nb_taps-1) of signed(11 downto 0);                
signal fir_reg                          : fir_reg_type:=(others=>(others=>'0'));                        
type taps_x_fir_reg_type                is array (0 to nb_taps-1) of signed(25 downto 0);                
signal taps_x_fir_reg                   : taps_x_fir_reg_type;                                           
                                                                                                         
type adder_tree_subtype                 is array (0 to nb_taps) of signed(63 downto 0);                  
type adder_tree_type                    is array (0 to nb_taps-1) of adder_tree_subtype;                 
signal adder_tree                       : adder_tree_type:=(others=>(others=>(others=>'0')));          
signal adder_tree_en                    : std_logic_vector(nb_taps-1 downto 0);                          
                                                                                                         
                                                                                                         
signal data_in_en_r1               : std_logic;                                                          
signal data_in_en_r2               : std_logic;                                                          
signal data_in_en_r3               : std_logic;                                                          
signal data_out_prepare            : std_logic_vector(11 downto 0);                                      
signal data_out_prepare_en         : std_logic;                                                          
                                                                                                         
begin                                                                                                    
                                                                                                         
                                                                                                         
                                                                                                         
    ------------------------------------------                                                           
    -- Fir implementation                                                                                
    ------------------------------------------                                                           
    process(clk)                                                                                         
    variable v_round : signed(1 downto 0);                                                               
    begin                                                                                                
                                                                                                         
        if rising_edge(clk) then                                                                         
                                                                                                         
            --shift registers                                                                            
            if data_in_en='1' then                                                                     
                fir_reg(0) <= signed(data_in);                                                           
                for I in 1 to nb_taps-1 loop                                                             
                       fir_reg(I) <= fir_reg(I-1);                                                       
                    end loop;                                                                            
            end if;                                                                                      
            data_in_en_r1 <= data_in_en;                                                                 
                                                                                                         
            --multiply                                                                                   
            for I in 0 to nb_taps-1 loop                                                                 
                taps_x_fir_reg(I) <= fir_reg(I) * taps(I); -- 12 + 14 = 26 bits                          
            end loop;                                                                                    
            data_in_en_r2 <= data_in_en_r1;                                                              
                                                                                                         
            --Pipe                                                                                       
            for I in 0 to nb_taps-1 loop                                                                 
                adder_tree(0)(I)         <= resize(taps_x_fir_reg(I),64);                                
            end loop;                                                                                    
            data_in_en_r3 <= data_in_en_r2;                                                              
                                                                                                         
            adder_tree(1)(0) <= adder_tree(0)(0) + adder_tree(0)(1); --27 bits 
            adder_tree(1)(1) <= adder_tree(0)(2) + adder_tree(0)(3); --27 bits 
            adder_tree(1)(2) <= adder_tree(0)(4) + adder_tree(0)(5); --27 bits 
            adder_tree(1)(3) <= adder_tree(0)(6) + adder_tree(0)(7); --27 bits 
            adder_tree(1)(4) <= adder_tree(0)(8) + adder_tree(0)(9); --27 bits 
            adder_tree(1)(5) <= adder_tree(0)(10) + adder_tree(0)(11); --27 bits 
            adder_tree(1)(6) <= adder_tree(0)(12) + adder_tree(0)(13); --27 bits 
            adder_tree(1)(7) <= adder_tree(0)(14) + adder_tree(0)(15); --27 bits 
            adder_tree(1)(8) <= adder_tree(0)(16) + adder_tree(0)(17); --27 bits 
            adder_tree(1)(9) <= adder_tree(0)(18) + adder_tree(0)(19); --27 bits 
            adder_tree(1)(10) <= adder_tree(0)(20) + adder_tree(0)(21); --27 bits 
            adder_tree(1)(11) <= adder_tree(0)(22) + adder_tree(0)(23); --27 bits 
            adder_tree(1)(12) <= adder_tree(0)(24) + adder_tree(0)(25); --27 bits 
            adder_tree(1)(13) <= adder_tree(0)(26) + adder_tree(0)(27); --27 bits 
            adder_tree(1)(14) <= adder_tree(0)(28) + adder_tree(0)(29); --27 bits 
            adder_tree(1)(15) <= adder_tree(0)(30) + adder_tree(0)(31); --27 bits 
            adder_tree(1)(16) <= adder_tree(0)(32) + adder_tree(0)(33); --27 bits 
            adder_tree(1)(17) <= adder_tree(0)(34) + adder_tree(0)(35); --27 bits 
            adder_tree(1)(18) <= adder_tree(0)(36) + adder_tree(0)(37); --27 bits 
            adder_tree(1)(19) <= adder_tree(0)(38) + adder_tree(0)(39); --27 bits 
            adder_tree(1)(20) <= adder_tree(0)(40) + adder_tree(0)(41); --27 bits 
            adder_tree(1)(21) <= adder_tree(0)(42) + adder_tree(0)(43); --27 bits 
            adder_tree(1)(22) <= adder_tree(0)(44) + adder_tree(0)(45); --27 bits 
            adder_tree(1)(23) <= adder_tree(0)(46) + adder_tree(0)(47); --27 bits 
            adder_tree(1)(24) <= adder_tree(0)(48) + adder_tree(0)(49); --27 bits 
            adder_tree(1)(25) <= adder_tree(0)(50) + adder_tree(0)(51); --27 bits 
            adder_tree(1)(26) <= adder_tree(0)(52) + adder_tree(0)(53); --27 bits 
            adder_tree(1)(27) <= adder_tree(0)(54) + adder_tree(0)(55); --27 bits 
            adder_tree(1)(28) <= adder_tree(0)(56) + adder_tree(0)(57); --27 bits 
            adder_tree(1)(29) <= adder_tree(0)(58) + adder_tree(0)(59); --27 bits 
            adder_tree(1)(30) <= adder_tree(0)(60) + adder_tree(0)(61); --27 bits 
            adder_tree(1)(31) <= adder_tree(0)(62) + adder_tree(0)(63); --27 bits 
            adder_tree(1)(32) <= adder_tree(0)(64) + adder_tree(0)(65); --27 bits 
            adder_tree(1)(33) <= adder_tree(0)(66) + adder_tree(0)(67); --27 bits 
            adder_tree(1)(34) <= adder_tree(0)(68) + adder_tree(0)(69); --27 bits 
            adder_tree(1)(35) <= adder_tree(0)(70) + adder_tree(0)(71); --27 bits 
            adder_tree(1)(36) <= adder_tree(0)(72) + adder_tree(0)(73); --27 bits 
            adder_tree(1)(37) <= adder_tree(0)(74) + adder_tree(0)(75); --27 bits 
            adder_tree(1)(38) <= adder_tree(0)(76) + adder_tree(0)(77); --27 bits 
            adder_tree(1)(39) <= adder_tree(0)(78) + adder_tree(0)(79); --27 bits 
            adder_tree(1)(40) <= adder_tree(0)(80) + adder_tree(0)(81); --27 bits 
            adder_tree(1)(41) <= adder_tree(0)(82) + adder_tree(0)(83); --27 bits 
            adder_tree(1)(42) <= adder_tree(0)(84) + adder_tree(0)(85); --27 bits 
            adder_tree(1)(43) <= adder_tree(0)(86) + adder_tree(0)(87); --27 bits 
            adder_tree(1)(44) <= adder_tree(0)(88) + adder_tree(0)(89); --27 bits 
            adder_tree(1)(45) <= adder_tree(0)(90) + adder_tree(0)(91); --27 bits 
            adder_tree(1)(46) <= adder_tree(0)(92) + adder_tree(0)(93); --27 bits 
            adder_tree(1)(47) <= adder_tree(0)(94) + adder_tree(0)(95); --27 bits 
            adder_tree(1)(48) <= adder_tree(0)(96) + adder_tree(0)(97); --27 bits 
            adder_tree(1)(49) <= adder_tree(0)(98) + adder_tree(0)(99); --27 bits 
            adder_tree(1)(50) <= adder_tree(0)(100) + adder_tree(0)(101); --27 bits 
            adder_tree(1)(51) <= adder_tree(0)(102) + adder_tree(0)(103); --27 bits 
            adder_tree(1)(52) <= adder_tree(0)(104) + adder_tree(0)(105); --27 bits 
            adder_tree(1)(53) <= adder_tree(0)(106) + adder_tree(0)(107); --27 bits 
            adder_tree(1)(54) <= adder_tree(0)(108) + adder_tree(0)(109); --27 bits 
            adder_tree(1)(55) <= adder_tree(0)(110) + adder_tree(0)(111); --27 bits 
            adder_tree(1)(56) <= adder_tree(0)(112) + adder_tree(0)(113); --27 bits 
            adder_tree(1)(57) <= adder_tree(0)(114) + adder_tree(0)(115); --27 bits 
            adder_tree(1)(58) <= adder_tree(0)(116) + adder_tree(0)(117); --27 bits 
            adder_tree(1)(59) <= adder_tree(0)(118) + adder_tree(0)(119); --27 bits 
            adder_tree(1)(60) <= adder_tree(0)(120) + adder_tree(0)(121); --27 bits 
            adder_tree(1)(61) <= adder_tree(0)(122) + adder_tree(0)(123); --27 bits 
            adder_tree(1)(62) <= adder_tree(0)(124) + adder_tree(0)(125); --27 bits 
            adder_tree(1)(63) <= adder_tree(0)(126) + adder_tree(0)(127); --27 bits 
            adder_tree(1)(64) <= adder_tree(0)(128) + adder_tree(0)(129); --27 bits 
            adder_tree(1)(65) <= adder_tree(0)(130) + adder_tree(0)(131); --27 bits 
            adder_tree(1)(66) <= adder_tree(0)(132) + adder_tree(0)(133); --27 bits 
            adder_tree(1)(67) <= adder_tree(0)(134) + adder_tree(0)(135); --27 bits 
            adder_tree(1)(68) <= adder_tree(0)(136) + adder_tree(0)(137); --27 bits 
            adder_tree(1)(69) <= adder_tree(0)(138) + adder_tree(0)(139); --27 bits 
            adder_tree(1)(70) <= adder_tree(0)(140) + adder_tree(0)(141); --27 bits 
            adder_tree(1)(71) <= adder_tree(0)(142) + adder_tree(0)(143); --27 bits 
            adder_tree(1)(72) <= adder_tree(0)(144) + adder_tree(0)(145); --27 bits 
            adder_tree(1)(73) <= adder_tree(0)(146) + adder_tree(0)(147); --27 bits 
            adder_tree(1)(74) <= adder_tree(0)(148) + adder_tree(0)(149); --27 bits 
            adder_tree(1)(75) <= adder_tree(0)(150) + adder_tree(0)(151); --27 bits 
            adder_tree(1)(76) <= adder_tree(0)(152) + adder_tree(0)(153); --27 bits 
            adder_tree(1)(77) <= adder_tree(0)(154) + adder_tree(0)(155); --27 bits 
            adder_tree(1)(78) <= adder_tree(0)(156) + adder_tree(0)(157); --27 bits 
            adder_tree(1)(79) <= adder_tree(0)(158) + adder_tree(0)(159); --27 bits 
            adder_tree(1)(80) <= adder_tree(0)(160) + adder_tree(0)(161); --27 bits 
            adder_tree(1)(81) <= adder_tree(0)(162) + adder_tree(0)(163); --27 bits 
            adder_tree(1)(82) <= adder_tree(0)(164) + adder_tree(0)(165); --27 bits 
            adder_tree(1)(83) <= adder_tree(0)(166) + adder_tree(0)(167); --27 bits 
            adder_tree(1)(84) <= adder_tree(0)(168) + adder_tree(0)(169); --27 bits 
            adder_tree(1)(85) <= adder_tree(0)(170) + adder_tree(0)(171); --27 bits 
            adder_tree(1)(86) <= adder_tree(0)(172) + adder_tree(0)(173); --27 bits 
            adder_tree(1)(87) <= adder_tree(0)(174) + adder_tree(0)(175); --27 bits 
            adder_tree(1)(88) <= adder_tree(0)(176) + adder_tree(0)(177); --27 bits 
            adder_tree(1)(89) <= adder_tree(0)(178) + adder_tree(0)(179); --27 bits 
            adder_tree(1)(90) <= adder_tree(0)(180) + adder_tree(0)(181); --27 bits 
            adder_tree(1)(91) <= adder_tree(0)(182) + adder_tree(0)(183); --27 bits 
            adder_tree(1)(92) <= adder_tree(0)(184) + adder_tree(0)(185); --27 bits 
            adder_tree(1)(93) <= adder_tree(0)(186) + adder_tree(0)(187); --27 bits 
            adder_tree(1)(94) <= adder_tree(0)(188) + adder_tree(0)(189); --27 bits 
            adder_tree(1)(95) <= adder_tree(0)(190) + adder_tree(0)(191); --27 bits 
            adder_tree(1)(96) <= adder_tree(0)(192) + adder_tree(0)(193); --27 bits 
            adder_tree(1)(97) <= adder_tree(0)(194) + adder_tree(0)(195); --27 bits 
            adder_tree(1)(98) <= adder_tree(0)(196) + adder_tree(0)(197); --27 bits 
            adder_tree(1)(99) <= adder_tree(0)(198) + adder_tree(0)(199); --27 bits 
            adder_tree(1)(100) <= adder_tree(0)(200) + adder_tree(0)(201); --27 bits 
            adder_tree(1)(101) <= adder_tree(0)(202) + adder_tree(0)(203); --27 bits 
            adder_tree(1)(102) <= adder_tree(0)(204) + adder_tree(0)(205); --27 bits 
            adder_tree(1)(103) <= adder_tree(0)(206) + adder_tree(0)(207); --27 bits 
            adder_tree(1)(104) <= adder_tree(0)(208) + adder_tree(0)(209); --27 bits 
            adder_tree(1)(105) <= adder_tree(0)(210) + adder_tree(0)(211); --27 bits 
            adder_tree(1)(106) <= adder_tree(0)(212) + adder_tree(0)(213); --27 bits 
            adder_tree(1)(107) <= adder_tree(0)(214) + adder_tree(0)(215); --27 bits 
            adder_tree(1)(108) <= adder_tree(0)(216) + adder_tree(0)(217); --27 bits 
            adder_tree(1)(109) <= adder_tree(0)(218) + adder_tree(0)(219); --27 bits 
            adder_tree(1)(110) <= adder_tree(0)(220) + adder_tree(0)(221); --27 bits 
            adder_tree(1)(111) <= adder_tree(0)(222) + adder_tree(0)(223); --27 bits 
            adder_tree(1)(112) <= adder_tree(0)(224) + adder_tree(0)(225); --27 bits 
            adder_tree(1)(113) <= adder_tree(0)(226) + adder_tree(0)(227); --27 bits 
            adder_tree(1)(114) <= adder_tree(0)(228) + adder_tree(0)(229); --27 bits 
            adder_tree(1)(115) <= adder_tree(0)(230) + adder_tree(0)(231); --27 bits 
            adder_tree(1)(116) <= adder_tree(0)(232) + adder_tree(0)(233); --27 bits 
            adder_tree(1)(117) <= adder_tree(0)(234) + adder_tree(0)(235); --27 bits 
            adder_tree(1)(118) <= adder_tree(0)(236) + adder_tree(0)(237); --27 bits 
            adder_tree(1)(119) <= adder_tree(0)(238) + adder_tree(0)(239); --27 bits 
            adder_tree(1)(120) <= adder_tree(0)(240) + adder_tree(0)(241); --27 bits 
            adder_tree(1)(121) <= adder_tree(0)(242) + adder_tree(0)(243); --27 bits 
            adder_tree(1)(122) <= adder_tree(0)(244) + adder_tree(0)(245); --27 bits 
            adder_tree(1)(123) <= adder_tree(0)(246) + adder_tree(0)(247); --27 bits 
            adder_tree(1)(124) <= adder_tree(0)(248) + adder_tree(0)(249); --27 bits 
            adder_tree(1)(125) <= adder_tree(0)(250) + adder_tree(0)(251); --27 bits 
            adder_tree(1)(126) <= adder_tree(0)(252) + adder_tree(0)(253); --27 bits 
            adder_tree(1)(127) <= adder_tree(0)(254) + adder_tree(0)(255); --27 bits 
            adder_tree(1)(128) <= adder_tree(0)(256) + adder_tree(0)(257); --27 bits 
            adder_tree(1)(129) <= adder_tree(0)(258) + adder_tree(0)(259); --27 bits 
            adder_tree(1)(130) <= adder_tree(0)(260) + adder_tree(0)(261); --27 bits 
            adder_tree(1)(131) <= adder_tree(0)(262) + adder_tree(0)(263); --27 bits 
            adder_tree(1)(132) <= adder_tree(0)(264) + adder_tree(0)(265); --27 bits 
            adder_tree(1)(133) <= adder_tree(0)(266) + adder_tree(0)(267); --27 bits 
            adder_tree(1)(134) <= adder_tree(0)(268) + adder_tree(0)(269); --27 bits 
            adder_tree(1)(135) <= adder_tree(0)(270) + adder_tree(0)(271); --27 bits 
            adder_tree(1)(136) <= adder_tree(0)(272) + adder_tree(0)(273); --27 bits 
            adder_tree(1)(137) <= adder_tree(0)(274) + adder_tree(0)(275); --27 bits 
            adder_tree(1)(138) <= adder_tree(0)(276) + adder_tree(0)(277); --27 bits 
            adder_tree(1)(139) <= adder_tree(0)(278) + adder_tree(0)(279); --27 bits 
            adder_tree(1)(140) <= adder_tree(0)(280) + adder_tree(0)(281); --27 bits 
            adder_tree(1)(141) <= adder_tree(0)(282) + adder_tree(0)(283); --27 bits 
            adder_tree(1)(142) <= adder_tree(0)(284) + adder_tree(0)(285); --27 bits 
            adder_tree(1)(143) <= adder_tree(0)(286) + adder_tree(0)(287); --27 bits 
            adder_tree(1)(144) <= adder_tree(0)(288) + adder_tree(0)(289); --27 bits 
            adder_tree(1)(145) <= adder_tree(0)(290) + adder_tree(0)(291); --27 bits 
            adder_tree(1)(146) <= adder_tree(0)(292) + adder_tree(0)(293); --27 bits 
            adder_tree(1)(147) <= adder_tree(0)(294) + adder_tree(0)(295); --27 bits 
            adder_tree(1)(148) <= adder_tree(0)(296) + adder_tree(0)(297); --27 bits 
            adder_tree(1)(149) <= adder_tree(0)(298) + adder_tree(0)(299); --27 bits 
            adder_tree(1)(150) <= adder_tree(0)(300) + adder_tree(0)(301); --27 bits 
            adder_tree(1)(151) <= adder_tree(0)(302) + adder_tree(0)(303); --27 bits 
            adder_tree(1)(152) <= adder_tree(0)(304) + adder_tree(0)(305); --27 bits 
            adder_tree(1)(153) <= adder_tree(0)(306) + adder_tree(0)(307); --27 bits 
            adder_tree(1)(154) <= adder_tree(0)(308) + adder_tree(0)(309); --27 bits 
            adder_tree(1)(155) <= adder_tree(0)(310) + adder_tree(0)(311); --27 bits 
            adder_tree(1)(156) <= adder_tree(0)(312) + adder_tree(0)(313); --27 bits 
            adder_tree(1)(157) <= adder_tree(0)(314) + adder_tree(0)(315); --27 bits 
            adder_tree(1)(158) <= adder_tree(0)(316) + adder_tree(0)(317); --27 bits 
            adder_tree(1)(159) <= adder_tree(0)(318) + adder_tree(0)(319); --27 bits 
            adder_tree(1)(160) <= adder_tree(0)(320) + adder_tree(0)(321); --27 bits 
            adder_tree(1)(161) <= adder_tree(0)(322) + adder_tree(0)(323); --27 bits 
            adder_tree(1)(162) <= adder_tree(0)(324) + adder_tree(0)(325); --27 bits 
            adder_tree(1)(163) <= adder_tree(0)(326) + adder_tree(0)(327); --27 bits 
            adder_tree(1)(164) <= adder_tree(0)(328) + adder_tree(0)(329); --27 bits 
            adder_tree(1)(165) <= adder_tree(0)(330) + adder_tree(0)(331); --27 bits 
            adder_tree(1)(166) <= adder_tree(0)(332) + adder_tree(0)(333); --27 bits 
            adder_tree(1)(167) <= adder_tree(0)(334) + adder_tree(0)(335); --27 bits 
            adder_tree(1)(168) <= adder_tree(0)(336) + adder_tree(0)(337); --27 bits 
            adder_tree(1)(169) <= adder_tree(0)(338) + adder_tree(0)(339); --27 bits 
            adder_tree(1)(170) <= adder_tree(0)(340) + adder_tree(0)(341); --27 bits 
            adder_tree(1)(171) <= adder_tree(0)(342) + adder_tree(0)(343); --27 bits 
            adder_tree(1)(172) <= adder_tree(0)(344) + adder_tree(0)(345); --27 bits 
            adder_tree(1)(173) <= adder_tree(0)(346) + adder_tree(0)(347); --27 bits 
            adder_tree(1)(174) <= adder_tree(0)(348) + adder_tree(0)(349); --27 bits 
            adder_tree(1)(175) <= adder_tree(0)(350) + adder_tree(0)(351); --27 bits 
            adder_tree(1)(176) <= adder_tree(0)(352) + adder_tree(0)(353); --27 bits 
            adder_tree(1)(177) <= adder_tree(0)(354) + adder_tree(0)(355); --27 bits 
            adder_tree(1)(178) <= adder_tree(0)(356) + adder_tree(0)(357); --27 bits 
            adder_tree(1)(179) <= adder_tree(0)(358) + adder_tree(0)(359); --27 bits 
            adder_tree(1)(180) <= adder_tree(0)(360) + adder_tree(0)(361); --27 bits 
            adder_tree(1)(181) <= adder_tree(0)(362) + adder_tree(0)(363); --27 bits 
            adder_tree(1)(182) <= adder_tree(0)(364) + adder_tree(0)(365); --27 bits 
            adder_tree(1)(183) <= adder_tree(0)(366) + adder_tree(0)(367); --27 bits 
            adder_tree(1)(184) <= adder_tree(0)(368) + adder_tree(0)(369); --27 bits 
            adder_tree(1)(185) <= adder_tree(0)(370) + adder_tree(0)(371); --27 bits 
            adder_tree(1)(186) <= adder_tree(0)(372) + adder_tree(0)(373); --27 bits 
            adder_tree(1)(187) <= adder_tree(0)(374) + adder_tree(0)(375); --27 bits 
            adder_tree(1)(188) <= adder_tree(0)(376) + adder_tree(0)(377); --27 bits 
            adder_tree(1)(189) <= adder_tree(0)(378) + adder_tree(0)(379); --27 bits 
            adder_tree(1)(190) <= adder_tree(0)(380) + adder_tree(0)(381); --27 bits 
            adder_tree(1)(191) <= adder_tree(0)(382) + adder_tree(0)(383); --27 bits 
            adder_tree(1)(192) <= adder_tree(0)(384) + adder_tree(0)(385); --27 bits 
            adder_tree(1)(193) <= adder_tree(0)(386) + adder_tree(0)(387); --27 bits 
            adder_tree(1)(194) <= adder_tree(0)(388) + adder_tree(0)(389); --27 bits 
            adder_tree(1)(195) <= adder_tree(0)(390) + adder_tree(0)(391); --27 bits 
            adder_tree(1)(196) <= adder_tree(0)(392) + adder_tree(0)(393); --27 bits 
            adder_tree(1)(197) <= adder_tree(0)(394) + adder_tree(0)(395); --27 bits 
            adder_tree(1)(198) <= adder_tree(0)(396) + adder_tree(0)(397); --27 bits 
            adder_tree(1)(199) <= adder_tree(0)(398) + adder_tree(0)(399); --27 bits 
            adder_tree(1)(200) <= adder_tree(0)(400) + adder_tree(0)(401); --27 bits 
            adder_tree(1)(201) <= adder_tree(0)(402) + adder_tree(0)(403); --27 bits 
            adder_tree(1)(202) <= adder_tree(0)(404) + adder_tree(0)(405); --27 bits 
            adder_tree(1)(203) <= adder_tree(0)(406) + adder_tree(0)(407); --27 bits 
            adder_tree(1)(204) <= adder_tree(0)(408) + adder_tree(0)(409); --27 bits 
            adder_tree(1)(205) <= adder_tree(0)(410) + adder_tree(0)(411); --27 bits 
            adder_tree(1)(206) <= adder_tree(0)(412) + adder_tree(0)(413); --27 bits 
            adder_tree(1)(207) <= adder_tree(0)(414) + adder_tree(0)(415); --27 bits 
            adder_tree(1)(208) <= adder_tree(0)(416) + adder_tree(0)(417); --27 bits 
            adder_tree(1)(209) <= adder_tree(0)(418) + adder_tree(0)(419); --27 bits 
            adder_tree(1)(210) <= adder_tree(0)(420) + adder_tree(0)(421); --27 bits 
            adder_tree(1)(211) <= adder_tree(0)(422) + adder_tree(0)(423); --27 bits 
            adder_tree(1)(212) <= adder_tree(0)(424) + adder_tree(0)(425); --27 bits 
            adder_tree(1)(213) <= adder_tree(0)(426) + adder_tree(0)(427); --27 bits 
            adder_tree(1)(214) <= adder_tree(0)(428) + adder_tree(0)(429); --27 bits 
            adder_tree(1)(215) <= adder_tree(0)(430) + adder_tree(0)(431); --27 bits 
            adder_tree(1)(216) <= adder_tree(0)(432) + adder_tree(0)(433); --27 bits 
            adder_tree(1)(217) <= adder_tree(0)(434) + adder_tree(0)(435); --27 bits 
            adder_tree(1)(218) <= adder_tree(0)(436) + adder_tree(0)(437); --27 bits 
            adder_tree(1)(219) <= adder_tree(0)(438) + adder_tree(0)(439); --27 bits 
            adder_tree(1)(220) <= adder_tree(0)(440) + adder_tree(0)(441); --27 bits 
            adder_tree(1)(221) <= adder_tree(0)(442) + adder_tree(0)(443); --27 bits 
            adder_tree(1)(222) <= adder_tree(0)(444) + adder_tree(0)(445); --27 bits 
            adder_tree(1)(223) <= adder_tree(0)(446) + adder_tree(0)(447); --27 bits 
            adder_tree(1)(224) <= adder_tree(0)(448) + adder_tree(0)(449); --27 bits 
            adder_tree(1)(225) <= adder_tree(0)(450) + adder_tree(0)(451); --27 bits 
            adder_tree(1)(226) <= adder_tree(0)(452) + adder_tree(0)(453); --27 bits 
            adder_tree(1)(227) <= adder_tree(0)(454) + adder_tree(0)(455); --27 bits 
            adder_tree(1)(228) <= adder_tree(0)(456) + adder_tree(0)(457); --27 bits 
            adder_tree(1)(229) <= adder_tree(0)(458) + adder_tree(0)(459); --27 bits 
            adder_tree(1)(230) <= adder_tree(0)(460) + adder_tree(0)(461); --27 bits 
            adder_tree(1)(231) <= adder_tree(0)(462) + adder_tree(0)(463); --27 bits 
            adder_tree(1)(232) <= adder_tree(0)(464) + adder_tree(0)(465); --27 bits 
            adder_tree(1)(233) <= adder_tree(0)(466) + adder_tree(0)(467); --27 bits 
            adder_tree(1)(234) <= adder_tree(0)(468) + adder_tree(0)(469); --27 bits 
            adder_tree(1)(235) <= adder_tree(0)(470) + adder_tree(0)(471); --27 bits 
            adder_tree(1)(236) <= adder_tree(0)(472) + adder_tree(0)(473); --27 bits 
            adder_tree(1)(237) <= adder_tree(0)(474) + adder_tree(0)(475); --27 bits 
            adder_tree(1)(238) <= adder_tree(0)(476) + adder_tree(0)(477); --27 bits 
            adder_tree(1)(239) <= adder_tree(0)(478) + adder_tree(0)(479); --27 bits 
            adder_tree(1)(240) <= adder_tree(0)(480) + adder_tree(0)(481); --27 bits 
            adder_tree(1)(241) <= adder_tree(0)(482) + adder_tree(0)(483); --27 bits 
            adder_tree(1)(242) <= adder_tree(0)(484) + adder_tree(0)(485); --27 bits 
            adder_tree(1)(243) <= adder_tree(0)(486) + adder_tree(0)(487); --27 bits 
            adder_tree(1)(244) <= adder_tree(0)(488) + adder_tree(0)(489); --27 bits 
            adder_tree(1)(245) <= adder_tree(0)(490) + adder_tree(0)(491); --27 bits 
            adder_tree(1)(246) <= adder_tree(0)(492) + adder_tree(0)(493); --27 bits 
            adder_tree(1)(247) <= adder_tree(0)(494) + adder_tree(0)(495); --27 bits 
            adder_tree(1)(248) <= adder_tree(0)(496) + adder_tree(0)(497); --27 bits 
            adder_tree(1)(249) <= adder_tree(0)(498) + adder_tree(0)(499); --27 bits 
            adder_tree(1)(250) <= adder_tree(0)(500) + adder_tree(0)(501); --27 bits 
            adder_tree(1)(251) <= adder_tree(0)(502) + adder_tree(0)(503); --27 bits 
            adder_tree(1)(252) <= adder_tree(0)(504) + adder_tree(0)(505); --27 bits 
            adder_tree(1)(253) <= adder_tree(0)(506) + adder_tree(0)(507); --27 bits 
            adder_tree(1)(254) <= adder_tree(0)(508) + adder_tree(0)(509); --27 bits 
            adder_tree(1)(255) <= adder_tree(0)(510) + adder_tree(0)(511); --27 bits 
            adder_tree(1)(256) <= adder_tree(0)(512) + adder_tree(0)(513); --27 bits 
            adder_tree(1)(257) <= adder_tree(0)(514) + adder_tree(0)(515); --27 bits 
            adder_tree(1)(258) <= adder_tree(0)(516) + adder_tree(0)(517); --27 bits 
            adder_tree(1)(259) <= adder_tree(0)(518) + adder_tree(0)(519); --27 bits 
            adder_tree(1)(260) <= adder_tree(0)(520) + adder_tree(0)(521); --27 bits 
            adder_tree(1)(261) <= adder_tree(0)(522) + adder_tree(0)(523); --27 bits 
            adder_tree(1)(262) <= adder_tree(0)(524) + adder_tree(0)(525); --27 bits 
            adder_tree(1)(263) <= adder_tree(0)(526) + adder_tree(0)(527); --27 bits 
            adder_tree(1)(264) <= adder_tree(0)(528) + adder_tree(0)(529); --27 bits 
            adder_tree(1)(265) <= adder_tree(0)(530) + adder_tree(0)(531); --27 bits 
            adder_tree(1)(266) <= adder_tree(0)(532) + adder_tree(0)(533); --27 bits 
            adder_tree(1)(267) <= adder_tree(0)(534) + adder_tree(0)(535); --27 bits 
            adder_tree(1)(268) <= adder_tree(0)(536) + adder_tree(0)(537); --27 bits 
            adder_tree(1)(269) <= adder_tree(0)(538) + adder_tree(0)(539); --27 bits 
            adder_tree(1)(270) <= adder_tree(0)(540) + adder_tree(0)(541); --27 bits 
            adder_tree(1)(271) <= adder_tree(0)(542) + adder_tree(0)(543); --27 bits 
            adder_tree(1)(272) <= adder_tree(0)(544) + adder_tree(0)(545); --27 bits 
            adder_tree(1)(273) <= adder_tree(0)(546) + adder_tree(0)(547); --27 bits 
            adder_tree(1)(274) <= adder_tree(0)(548) + adder_tree(0)(549); --27 bits 
            adder_tree(1)(275) <= adder_tree(0)(550) + adder_tree(0)(551); --27 bits 
            adder_tree(1)(276) <= adder_tree(0)(552) + adder_tree(0)(553); --27 bits 
            adder_tree(1)(277) <= adder_tree(0)(554) + adder_tree(0)(555); --27 bits 
            adder_tree(1)(278) <= adder_tree(0)(556) + adder_tree(0)(557); --27 bits 
            adder_tree(1)(279) <= adder_tree(0)(558) + adder_tree(0)(559); --27 bits 
            adder_tree(1)(280) <= adder_tree(0)(560) + adder_tree(0)(561); --27 bits 
            adder_tree(1)(281) <= adder_tree(0)(562) + adder_tree(0)(563); --27 bits 
            adder_tree(1)(282) <= adder_tree(0)(564) + adder_tree(0)(565); --27 bits 
            adder_tree(1)(283) <= adder_tree(0)(566) + adder_tree(0)(567); --27 bits 
            adder_tree(1)(284) <= adder_tree(0)(568) + adder_tree(0)(569); --27 bits 
            adder_tree(1)(285) <= adder_tree(0)(570) + adder_tree(0)(571); --27 bits 
            adder_tree(1)(286) <= adder_tree(0)(572) + adder_tree(0)(573); --27 bits 
            adder_tree(1)(287) <= adder_tree(0)(574) + adder_tree(0)(575); --27 bits 
            adder_tree(1)(288) <= adder_tree(0)(576) + adder_tree(0)(577); --27 bits 
            adder_tree(1)(289) <= adder_tree(0)(578) + adder_tree(0)(579); --27 bits 
            adder_tree(1)(290) <= adder_tree(0)(580) + adder_tree(0)(581); --27 bits 
            adder_tree(1)(291) <= adder_tree(0)(582) + adder_tree(0)(583); --27 bits 
            adder_tree(1)(292) <= adder_tree(0)(584) + adder_tree(0)(585); --27 bits 
            adder_tree(1)(293) <= adder_tree(0)(586) + adder_tree(0)(587); --27 bits 
            adder_tree(1)(294) <= adder_tree(0)(588) + adder_tree(0)(589); --27 bits 
            adder_tree(1)(295) <= adder_tree(0)(590) + adder_tree(0)(591); --27 bits 
            adder_tree(1)(296) <= adder_tree(0)(592) + adder_tree(0)(593); --27 bits 
            adder_tree(1)(297) <= adder_tree(0)(594) + adder_tree(0)(595); --27 bits 
            adder_tree(1)(298) <= adder_tree(0)(596) + adder_tree(0)(597); --27 bits 
            adder_tree(1)(299) <= adder_tree(0)(598) + adder_tree(0)(599); --27 bits 
            adder_tree(1)(300) <= adder_tree(0)(600) + adder_tree(0)(601); --27 bits 
            adder_tree(1)(301) <= adder_tree(0)(602) + adder_tree(0)(603); --27 bits 
            adder_tree(1)(302) <= adder_tree(0)(604) + adder_tree(0)(605); --27 bits 
            adder_tree(1)(303) <= adder_tree(0)(606) + adder_tree(0)(607); --27 bits 
            adder_tree(1)(304) <= adder_tree(0)(608) + adder_tree(0)(609); --27 bits 
            adder_tree(1)(305) <= adder_tree(0)(610) + adder_tree(0)(611); --27 bits 
            adder_tree(1)(306) <= adder_tree(0)(612) + adder_tree(0)(613); --27 bits 
            adder_tree(1)(307) <= adder_tree(0)(614) + adder_tree(0)(615); --27 bits 
            adder_tree(1)(308) <= adder_tree(0)(616) + adder_tree(0)(617); --27 bits 
            adder_tree(1)(309) <= adder_tree(0)(618) + adder_tree(0)(619); --27 bits 
            adder_tree(1)(310) <= adder_tree(0)(620) + adder_tree(0)(621); --27 bits 
            adder_tree(1)(311) <= adder_tree(0)(622) + adder_tree(0)(623); --27 bits 
            adder_tree(1)(312) <= adder_tree(0)(624) + adder_tree(0)(625); --27 bits 
            adder_tree(1)(313) <= adder_tree(0)(626) + adder_tree(0)(627); --27 bits 
            adder_tree(1)(314) <= adder_tree(0)(628) + adder_tree(0)(629); --27 bits 
            adder_tree(1)(315) <= adder_tree(0)(630) + adder_tree(0)(631); --27 bits 
            adder_tree(1)(316) <= adder_tree(0)(632) + adder_tree(0)(633); --27 bits 
            adder_tree(1)(317) <= adder_tree(0)(634) + adder_tree(0)(635); --27 bits 
            adder_tree(1)(318) <= adder_tree(0)(636) + adder_tree(0)(637); --27 bits 
            adder_tree(1)(319) <= adder_tree(0)(638) + adder_tree(0)(639); --27 bits 
            adder_tree(1)(320) <= adder_tree(0)(640) + adder_tree(0)(641); --27 bits 
            adder_tree(1)(321) <= adder_tree(0)(642) + adder_tree(0)(643); --27 bits 
            adder_tree(1)(322) <= adder_tree(0)(644) + adder_tree(0)(645); --27 bits 
            adder_tree(1)(323) <= adder_tree(0)(646) + adder_tree(0)(647); --27 bits 
            adder_tree(1)(324) <= adder_tree(0)(648) + adder_tree(0)(649); --27 bits 
            adder_tree(1)(325) <= adder_tree(0)(650) + adder_tree(0)(651); --27 bits 
            adder_tree(1)(326) <= adder_tree(0)(652) + adder_tree(0)(653); --27 bits 
            adder_tree(1)(327) <= adder_tree(0)(654) + adder_tree(0)(655); --27 bits 
            adder_tree(1)(328) <= adder_tree(0)(656) + adder_tree(0)(657); --27 bits 
            adder_tree(1)(329) <= adder_tree(0)(658) + adder_tree(0)(659); --27 bits 
            adder_tree(1)(330) <= adder_tree(0)(660) + adder_tree(0)(661); --27 bits 
            adder_tree(1)(331) <= adder_tree(0)(662) + adder_tree(0)(663); --27 bits 
            adder_tree(1)(332) <= adder_tree(0)(664) + adder_tree(0)(665); --27 bits 
            adder_tree(1)(333) <= adder_tree(0)(666) + adder_tree(0)(667); --27 bits 
            adder_tree(1)(334) <= adder_tree(0)(668) + adder_tree(0)(669); --27 bits 
            adder_tree(1)(335) <= adder_tree(0)(670) + adder_tree(0)(671); --27 bits 
            adder_tree(1)(336) <= adder_tree(0)(672) + adder_tree(0)(673); --27 bits 
            adder_tree(1)(337) <= adder_tree(0)(674) + adder_tree(0)(675); --27 bits 
            adder_tree(1)(338) <= adder_tree(0)(676) + adder_tree(0)(677); --27 bits 
            adder_tree(1)(339) <= adder_tree(0)(678) + adder_tree(0)(679); --27 bits 
            adder_tree(1)(340) <= adder_tree(0)(680) + adder_tree(0)(681); --27 bits 
            adder_tree(1)(341) <= adder_tree(0)(682) + adder_tree(0)(683); --27 bits 
            adder_tree(1)(342) <= adder_tree(0)(684) + adder_tree(0)(685); --27 bits 
            adder_tree(1)(343) <= adder_tree(0)(686) + adder_tree(0)(687); --27 bits 
            adder_tree(1)(344) <= adder_tree(0)(688) + adder_tree(0)(689); --27 bits 
            adder_tree(1)(345) <= adder_tree(0)(690) + adder_tree(0)(691); --27 bits 
            adder_tree(1)(346) <= adder_tree(0)(692) + adder_tree(0)(693); --27 bits 
            adder_tree(1)(347) <= adder_tree(0)(694) + adder_tree(0)(695); --27 bits 
            adder_tree(1)(348) <= adder_tree(0)(696) + adder_tree(0)(697); --27 bits 
            adder_tree(1)(349) <= adder_tree(0)(698) + adder_tree(0)(699); --27 bits 
            adder_tree(1)(350) <= adder_tree(0)(700) + adder_tree(0)(701); --27 bits 
            adder_tree(1)(351) <= adder_tree(0)(702) + adder_tree(0)(703); --27 bits 
            adder_tree(1)(352) <= adder_tree(0)(704) + adder_tree(0)(705); --27 bits 
            adder_tree(1)(353) <= adder_tree(0)(706) + adder_tree(0)(707); --27 bits 
            adder_tree(1)(354) <= adder_tree(0)(708) + adder_tree(0)(709); --27 bits 
            adder_tree(1)(355) <= adder_tree(0)(710) + adder_tree(0)(711); --27 bits 
            adder_tree(1)(356) <= adder_tree(0)(712) + adder_tree(0)(713); --27 bits 
            adder_tree(1)(357) <= adder_tree(0)(714) + adder_tree(0)(715); --27 bits 
            adder_tree(1)(358) <= adder_tree(0)(716) + adder_tree(0)(717); --27 bits 
            adder_tree(1)(359) <= adder_tree(0)(718) + adder_tree(0)(719); --27 bits 
            adder_tree(1)(360) <= adder_tree(0)(720) + adder_tree(0)(721); --27 bits 
            adder_tree(1)(361) <= adder_tree(0)(722) + adder_tree(0)(723); --27 bits 
            adder_tree(1)(362) <= adder_tree(0)(724) + adder_tree(0)(725); --27 bits 
            adder_tree(1)(363) <= adder_tree(0)(726) + adder_tree(0)(727); --27 bits 
            adder_tree(1)(364) <= adder_tree(0)(728) + adder_tree(0)(729); --27 bits 
            adder_tree(1)(365) <= adder_tree(0)(730) + adder_tree(0)(731); --27 bits 
            adder_tree(1)(366) <= adder_tree(0)(732) + adder_tree(0)(733); --27 bits 
            adder_tree(1)(367) <= adder_tree(0)(734) + adder_tree(0)(735); --27 bits 
            adder_tree(1)(368) <= adder_tree(0)(736) + adder_tree(0)(737); --27 bits 
            adder_tree(1)(369) <= adder_tree(0)(738) + adder_tree(0)(739); --27 bits 
            adder_tree(1)(370) <= adder_tree(0)(740) + adder_tree(0)(741); --27 bits 
            adder_tree(1)(371) <= adder_tree(0)(742) + adder_tree(0)(743); --27 bits 
            adder_tree(1)(372) <= adder_tree(0)(744) + adder_tree(0)(745); --27 bits 
            adder_tree(1)(373) <= adder_tree(0)(746) + adder_tree(0)(747); --27 bits 
            adder_tree(1)(374) <= adder_tree(0)(748) + adder_tree(0)(749); --27 bits 
            adder_tree(1)(375) <= adder_tree(0)(750) + adder_tree(0)(751); --27 bits 
            adder_tree(1)(376) <= adder_tree(0)(752) + adder_tree(0)(753); --27 bits 
            adder_tree(1)(377) <= adder_tree(0)(754) + adder_tree(0)(755); --27 bits 
            adder_tree(1)(378) <= adder_tree(0)(756) + adder_tree(0)(757); --27 bits 
            adder_tree(1)(379) <= adder_tree(0)(758) + adder_tree(0)(759); --27 bits 
            adder_tree(1)(380) <= adder_tree(0)(760) + adder_tree(0)(761); --27 bits 
            adder_tree(1)(381) <= adder_tree(0)(762) + adder_tree(0)(763); --27 bits 
            adder_tree(1)(382) <= adder_tree(0)(764) + adder_tree(0)(765); --27 bits 
            adder_tree(1)(383) <= adder_tree(0)(766) + adder_tree(0)(767); --27 bits 
            adder_tree(1)(384) <= adder_tree(0)(768) + adder_tree(0)(769); --27 bits 
            adder_tree(1)(385) <= adder_tree(0)(770) + adder_tree(0)(771); --27 bits 
            adder_tree(1)(386) <= adder_tree(0)(772) + adder_tree(0)(773); --27 bits 
            adder_tree(1)(387) <= adder_tree(0)(774) + adder_tree(0)(775); --27 bits 
            adder_tree(1)(388) <= adder_tree(0)(776) + adder_tree(0)(777); --27 bits 
            adder_tree(1)(389) <= adder_tree(0)(778) + adder_tree(0)(779); --27 bits 
            adder_tree(1)(390) <= adder_tree(0)(780) + adder_tree(0)(781); --27 bits 
            adder_tree(1)(391) <= adder_tree(0)(782) + adder_tree(0)(783); --27 bits 
            adder_tree(1)(392) <= adder_tree(0)(784) + adder_tree(0)(785); --27 bits 
            adder_tree(1)(393) <= adder_tree(0)(786) + adder_tree(0)(787); --27 bits 
            adder_tree(1)(394) <= adder_tree(0)(788) + adder_tree(0)(789); --27 bits 
            adder_tree(1)(395) <= adder_tree(0)(790) + adder_tree(0)(791); --27 bits 
            adder_tree(1)(396) <= adder_tree(0)(792) + adder_tree(0)(793); --27 bits 
            adder_tree(1)(397) <= adder_tree(0)(794) + adder_tree(0)(795); --27 bits 
            adder_tree(1)(398) <= adder_tree(0)(796) + adder_tree(0)(797); --27 bits 
            adder_tree(1)(399) <= adder_tree(0)(798) + adder_tree(0)(799); --27 bits 
            adder_tree(1)(400) <= adder_tree(0)(800) + adder_tree(0)(801); --27 bits 
            adder_tree(1)(401) <= adder_tree(0)(802) + adder_tree(0)(803); --27 bits 
            adder_tree(1)(402) <= adder_tree(0)(804) + adder_tree(0)(805); --27 bits 
            adder_tree(1)(403) <= adder_tree(0)(806) + adder_tree(0)(807); --27 bits 
            adder_tree(1)(404) <= adder_tree(0)(808) + adder_tree(0)(809); --27 bits 
            adder_tree(1)(405) <= adder_tree(0)(810) + adder_tree(0)(811); --27 bits 
            adder_tree(1)(406) <= adder_tree(0)(812) + adder_tree(0)(813); --27 bits 
            adder_tree(1)(407) <= adder_tree(0)(814) + adder_tree(0)(815); --27 bits 
            adder_tree(1)(408) <= adder_tree(0)(816) + adder_tree(0)(817); --27 bits 
            adder_tree(1)(409) <= adder_tree(0)(818) + adder_tree(0)(819); --27 bits 
            adder_tree(1)(410) <= adder_tree(0)(820) + adder_tree(0)(821); --27 bits 
            adder_tree(1)(411) <= adder_tree(0)(822) + adder_tree(0)(823); --27 bits 
            adder_tree(1)(412) <= adder_tree(0)(824) + adder_tree(0)(825); --27 bits 
            adder_tree(1)(413) <= adder_tree(0)(826) + adder_tree(0)(827); --27 bits 
            adder_tree(1)(414) <= adder_tree(0)(828) + adder_tree(0)(829); --27 bits 
            adder_tree(1)(415) <= adder_tree(0)(830) + adder_tree(0)(831); --27 bits 
            adder_tree(1)(416) <= adder_tree(0)(832) + adder_tree(0)(833); --27 bits 
            adder_tree(1)(417) <= adder_tree(0)(834) + adder_tree(0)(835); --27 bits 
            adder_tree(1)(418) <= adder_tree(0)(836) + adder_tree(0)(837); --27 bits 
            adder_tree(1)(419) <= adder_tree(0)(838) + adder_tree(0)(839); --27 bits 
            adder_tree(1)(420) <= adder_tree(0)(840) + adder_tree(0)(841); --27 bits 
            adder_tree(1)(421) <= adder_tree(0)(842) + adder_tree(0)(843); --27 bits 
            adder_tree(1)(422) <= adder_tree(0)(844) + adder_tree(0)(845); --27 bits 
            adder_tree(1)(423) <= adder_tree(0)(846) + adder_tree(0)(847); --27 bits 
            adder_tree(1)(424) <= adder_tree(0)(848) + adder_tree(0)(849); --27 bits 
            adder_tree(1)(425) <= adder_tree(0)(850) + adder_tree(0)(851); --27 bits 
            adder_tree(1)(426) <= adder_tree(0)(852) + adder_tree(0)(853); --27 bits 
            adder_tree(1)(427) <= adder_tree(0)(854) + adder_tree(0)(855); --27 bits 
            adder_tree(1)(428) <= adder_tree(0)(856) + adder_tree(0)(857); --27 bits 
            adder_tree(1)(429) <= adder_tree(0)(858) + adder_tree(0)(859); --27 bits 
            adder_tree(1)(430) <= adder_tree(0)(860) + adder_tree(0)(861); --27 bits 
            adder_tree(1)(431) <= adder_tree(0)(862) + adder_tree(0)(863); --27 bits 
            adder_tree(1)(432) <= adder_tree(0)(864) + adder_tree(0)(865); --27 bits 
            adder_tree(1)(433) <= adder_tree(0)(866) + adder_tree(0)(867); --27 bits 
            adder_tree(1)(434) <= adder_tree(0)(868) + adder_tree(0)(869); --27 bits 
            adder_tree(1)(435) <= adder_tree(0)(870) + adder_tree(0)(871); --27 bits 
            adder_tree(1)(436) <= adder_tree(0)(872) + adder_tree(0)(873); --27 bits 
            adder_tree(1)(437) <= adder_tree(0)(874) + adder_tree(0)(875); --27 bits 
            adder_tree(1)(438) <= adder_tree(0)(876) + adder_tree(0)(877); --27 bits 
            adder_tree(1)(439) <= adder_tree(0)(878) + adder_tree(0)(879); --27 bits 
            adder_tree(1)(440) <= adder_tree(0)(880) + adder_tree(0)(881); --27 bits 
            adder_tree(1)(441) <= adder_tree(0)(882) + adder_tree(0)(883); --27 bits 
            adder_tree(1)(442) <= adder_tree(0)(884) + adder_tree(0)(885); --27 bits 
            adder_tree(1)(443) <= adder_tree(0)(886) + adder_tree(0)(887); --27 bits 
            adder_tree(1)(444) <= adder_tree(0)(888) + adder_tree(0)(889); --27 bits 
            adder_tree(1)(445) <= adder_tree(0)(890) + adder_tree(0)(891); --27 bits 
            adder_tree(1)(446) <= adder_tree(0)(892) + adder_tree(0)(893); --27 bits 
            adder_tree(1)(447) <= adder_tree(0)(894) + adder_tree(0)(895); --27 bits 
            adder_tree(1)(448) <= adder_tree(0)(896) + adder_tree(0)(897); --27 bits 
            adder_tree(1)(449) <= adder_tree(0)(898) + adder_tree(0)(899); --27 bits 
            adder_tree(1)(450) <= adder_tree(0)(900) + adder_tree(0)(901); --27 bits 
            adder_tree(1)(451) <= adder_tree(0)(902) + adder_tree(0)(903); --27 bits 
            adder_tree(1)(452) <= adder_tree(0)(904) + adder_tree(0)(905); --27 bits 
            adder_tree(1)(453) <= adder_tree(0)(906) + adder_tree(0)(907); --27 bits 
            adder_tree(1)(454) <= adder_tree(0)(908) + adder_tree(0)(909); --27 bits 
            adder_tree(1)(455) <= adder_tree(0)(910) + adder_tree(0)(911); --27 bits 
            adder_tree(1)(456) <= adder_tree(0)(912) + adder_tree(0)(913); --27 bits 
            adder_tree(1)(457) <= adder_tree(0)(914) + adder_tree(0)(915); --27 bits 
            adder_tree(1)(458) <= adder_tree(0)(916) + adder_tree(0)(917); --27 bits 
            adder_tree(1)(459) <= adder_tree(0)(918) + adder_tree(0)(919); --27 bits 
            adder_tree(1)(460) <= adder_tree(0)(920) + adder_tree(0)(921); --27 bits 
            adder_tree(1)(461) <= adder_tree(0)(922) + adder_tree(0)(923); --27 bits 
            adder_tree(1)(462) <= adder_tree(0)(924) + adder_tree(0)(925); --27 bits 
            adder_tree(1)(463) <= adder_tree(0)(926) + adder_tree(0)(927); --27 bits 
            adder_tree(1)(464) <= adder_tree(0)(928) + adder_tree(0)(929); --27 bits 
            adder_tree(1)(465) <= adder_tree(0)(930) + adder_tree(0)(931); --27 bits 
            adder_tree(1)(466) <= adder_tree(0)(932) + adder_tree(0)(933); --27 bits 
            adder_tree(1)(467) <= adder_tree(0)(934) + adder_tree(0)(935); --27 bits 
            adder_tree(1)(468) <= adder_tree(0)(936) + adder_tree(0)(937); --27 bits 
            adder_tree(1)(469) <= adder_tree(0)(938) + adder_tree(0)(939); --27 bits 
            adder_tree(1)(470) <= adder_tree(0)(940) + adder_tree(0)(941); --27 bits 
            adder_tree(1)(471) <= adder_tree(0)(942) + adder_tree(0)(943); --27 bits 
            adder_tree(1)(472) <= adder_tree(0)(944) + adder_tree(0)(945); --27 bits 
            adder_tree(1)(473) <= adder_tree(0)(946) + adder_tree(0)(947); --27 bits 
            adder_tree(1)(474) <= adder_tree(0)(948) + adder_tree(0)(949); --27 bits 
            adder_tree(1)(475) <= adder_tree(0)(950) + adder_tree(0)(951); --27 bits 
            adder_tree(1)(476) <= adder_tree(0)(952) + adder_tree(0)(953); --27 bits 
            adder_tree(1)(477) <= adder_tree(0)(954) + adder_tree(0)(955); --27 bits 
            adder_tree(1)(478) <= adder_tree(0)(956) + adder_tree(0)(957); --27 bits 
            adder_tree(1)(479) <= adder_tree(0)(958) + adder_tree(0)(959); --27 bits 
            adder_tree(1)(480) <= adder_tree(0)(960) + adder_tree(0)(961); --27 bits 
            adder_tree(1)(481) <= adder_tree(0)(962) + adder_tree(0)(963); --27 bits 
            adder_tree(1)(482) <= adder_tree(0)(964) + adder_tree(0)(965); --27 bits 
            adder_tree(1)(483) <= adder_tree(0)(966) + adder_tree(0)(967); --27 bits 
            adder_tree(1)(484) <= adder_tree(0)(968) + adder_tree(0)(969); --27 bits 
            adder_tree(1)(485) <= adder_tree(0)(970) + adder_tree(0)(971); --27 bits 
            adder_tree(1)(486) <= adder_tree(0)(972) + adder_tree(0)(973); --27 bits 
            adder_tree(1)(487) <= adder_tree(0)(974) + adder_tree(0)(975); --27 bits 
            adder_tree(1)(488) <= adder_tree(0)(976) + adder_tree(0)(977); --27 bits 
            adder_tree(1)(489) <= adder_tree(0)(978) + adder_tree(0)(979); --27 bits 
            adder_tree(1)(490) <= adder_tree(0)(980) + adder_tree(0)(981); --27 bits 
            adder_tree(1)(491) <= adder_tree(0)(982) + adder_tree(0)(983); --27 bits 
            adder_tree(1)(492) <= adder_tree(0)(984) + adder_tree(0)(985); --27 bits 
            adder_tree(1)(493) <= adder_tree(0)(986) + adder_tree(0)(987); --27 bits 
            adder_tree(1)(494) <= adder_tree(0)(988) + adder_tree(0)(989); --27 bits 
            adder_tree(1)(495) <= adder_tree(0)(990) + adder_tree(0)(991); --27 bits 
            adder_tree(1)(496) <= adder_tree(0)(992) + adder_tree(0)(993); --27 bits 
            adder_tree(1)(497) <= adder_tree(0)(994) + adder_tree(0)(995); --27 bits 
            adder_tree(1)(498) <= adder_tree(0)(996) + adder_tree(0)(997); --27 bits 
            adder_tree(1)(499) <= adder_tree(0)(998) + adder_tree(0)(999); --27 bits 
            adder_tree(1)(500) <= adder_tree(0)(1000) + adder_tree(0)(1001); --27 bits 
            adder_tree(1)(501) <= adder_tree(0)(1002) + adder_tree(0)(1003); --27 bits 
            adder_tree(1)(502) <= adder_tree(0)(1004) + adder_tree(0)(1005); --27 bits 
            adder_tree(1)(503) <= adder_tree(0)(1006) + adder_tree(0)(1007); --27 bits 
            adder_tree(1)(504) <= adder_tree(0)(1008) + adder_tree(0)(1009); --27 bits 
            adder_tree(1)(505) <= adder_tree(0)(1010) + adder_tree(0)(1011); --27 bits 
            adder_tree(1)(506) <= adder_tree(0)(1012) + adder_tree(0)(1013); --27 bits 
            adder_tree(1)(507) <= adder_tree(0)(1014) + adder_tree(0)(1015); --27 bits 
            adder_tree(1)(508) <= adder_tree(0)(1016) + adder_tree(0)(1017); --27 bits 
            adder_tree(1)(509) <= adder_tree(0)(1018) + adder_tree(0)(1019); --27 bits 
            adder_tree(1)(510) <= adder_tree(0)(1020) + adder_tree(0)(1021); --27 bits 
            adder_tree(1)(511) <= adder_tree(0)(1022) + adder_tree(0)(1023); --27 bits 
            adder_tree(1)(512) <= adder_tree(0)(1024) + adder_tree(0)(1025); --27 bits 
            adder_tree(1)(513) <= adder_tree(0)(1026) + adder_tree(0)(1027); --27 bits 
            adder_tree(1)(514) <= adder_tree(0)(1028) + adder_tree(0)(1029); --27 bits 
            adder_tree(1)(515) <= adder_tree(0)(1030) + adder_tree(0)(1031); --27 bits 
            adder_tree(1)(516) <= adder_tree(0)(1032) + adder_tree(0)(1033); --27 bits 
            adder_tree(1)(517) <= adder_tree(0)(1034) + adder_tree(0)(1035); --27 bits 
            adder_tree(1)(518) <= adder_tree(0)(1036) + adder_tree(0)(1037); --27 bits 
            adder_tree(1)(519) <= adder_tree(0)(1038) + adder_tree(0)(1039); --27 bits 
            adder_tree(1)(520) <= adder_tree(0)(1040) + adder_tree(0)(1041); --27 bits 
            adder_tree(1)(521) <= adder_tree(0)(1042) + adder_tree(0)(1043); --27 bits 
            adder_tree(1)(522) <= adder_tree(0)(1044) + adder_tree(0)(1045); --27 bits 
            adder_tree(1)(523) <= adder_tree(0)(1046) + adder_tree(0)(1047); --27 bits 
            adder_tree(1)(524) <= adder_tree(0)(1048) + adder_tree(0)(1049); --27 bits 
            adder_tree(1)(525) <= adder_tree(0)(1050) + adder_tree(0)(1051); --27 bits 
            adder_tree(1)(526) <= adder_tree(0)(1052) + adder_tree(0)(1053); --27 bits 
            adder_tree(1)(527) <= adder_tree(0)(1054) + adder_tree(0)(1055); --27 bits 
            adder_tree(1)(528) <= adder_tree(0)(1056) + adder_tree(0)(1057); --27 bits 
            adder_tree(1)(529) <= adder_tree(0)(1058) + adder_tree(0)(1059); --27 bits 
            adder_tree(1)(530) <= adder_tree(0)(1060) + adder_tree(0)(1061); --27 bits 
            adder_tree(1)(531) <= adder_tree(0)(1062) + adder_tree(0)(1063); --27 bits 
            adder_tree(1)(532) <= adder_tree(0)(1064) + adder_tree(0)(1065); --27 bits 
            adder_tree(1)(533) <= adder_tree(0)(1066) + adder_tree(0)(1067); --27 bits 
            adder_tree(1)(534) <= adder_tree(0)(1068) + adder_tree(0)(1069); --27 bits 
            adder_tree(1)(535) <= adder_tree(0)(1070) + adder_tree(0)(1071); --27 bits 
            adder_tree(1)(536) <= adder_tree(0)(1072) + adder_tree(0)(1073); --27 bits 
            adder_tree(1)(537) <= adder_tree(0)(1074) + adder_tree(0)(1075); --27 bits 
            adder_tree(1)(538) <= adder_tree(0)(1076) + adder_tree(0)(1077); --27 bits 
            adder_tree(1)(539) <= adder_tree(0)(1078) + adder_tree(0)(1079); --27 bits 
            adder_tree(1)(540) <= adder_tree(0)(1080) + adder_tree(0)(1081); --27 bits 
            adder_tree(1)(541) <= adder_tree(0)(1082) + adder_tree(0)(1083); --27 bits 
            adder_tree(1)(542) <= adder_tree(0)(1084) + adder_tree(0)(1085); --27 bits 
            adder_tree(1)(543) <= adder_tree(0)(1086) + adder_tree(0)(1087); --27 bits 
            adder_tree(1)(544) <= adder_tree(0)(1088) + adder_tree(0)(1089); --27 bits 
            adder_tree(1)(545) <= adder_tree(0)(1090) + adder_tree(0)(1091); --27 bits 
            adder_tree(1)(546) <= adder_tree(0)(1092) + adder_tree(0)(1093); --27 bits 
            adder_tree(1)(547) <= adder_tree(0)(1094) + adder_tree(0)(1095); --27 bits 
            adder_tree(1)(548) <= adder_tree(0)(1096) + adder_tree(0)(1097); --27 bits 
            adder_tree(1)(549) <= adder_tree(0)(1098) + adder_tree(0)(1099); --27 bits 
            adder_tree(1)(550) <= adder_tree(0)(1100) + adder_tree(0)(1101); --27 bits 
            adder_tree(1)(551) <= adder_tree(0)(1102) + adder_tree(0)(1103); --27 bits 
            adder_tree(1)(552) <= adder_tree(0)(1104) + adder_tree(0)(1105); --27 bits 
            adder_tree(1)(553) <= adder_tree(0)(1106) + adder_tree(0)(1107); --27 bits 
            adder_tree(1)(554) <= adder_tree(0)(1108) + adder_tree(0)(1109); --27 bits 
            adder_tree(1)(555) <= adder_tree(0)(1110) + adder_tree(0)(1111); --27 bits 
            adder_tree(1)(556) <= adder_tree(0)(1112) + adder_tree(0)(1113); --27 bits 
            adder_tree(1)(557) <= adder_tree(0)(1114) + adder_tree(0)(1115); --27 bits 
            adder_tree(1)(558) <= adder_tree(0)(1116) + adder_tree(0)(1117); --27 bits 
            adder_tree(1)(559) <= adder_tree(0)(1118) + adder_tree(0)(1119); --27 bits 
            adder_tree(1)(560) <= adder_tree(0)(1120) + adder_tree(0)(1121); --27 bits 
            adder_tree(1)(561) <= adder_tree(0)(1122) + adder_tree(0)(1123); --27 bits 
            adder_tree(1)(562) <= adder_tree(0)(1124) + adder_tree(0)(1125); --27 bits 
            adder_tree(1)(563) <= adder_tree(0)(1126) + adder_tree(0)(1127); --27 bits 
            adder_tree(1)(564) <= adder_tree(0)(1128) + adder_tree(0)(1129); --27 bits 
            adder_tree(1)(565) <= adder_tree(0)(1130) + adder_tree(0)(1131); --27 bits 
            adder_tree(1)(566) <= adder_tree(0)(1132) + adder_tree(0)(1133); --27 bits 
            adder_tree(1)(567) <= adder_tree(0)(1134) + adder_tree(0)(1135); --27 bits 
            adder_tree(1)(568) <= adder_tree(0)(1136) + adder_tree(0)(1137); --27 bits 
            adder_tree(1)(569) <= adder_tree(0)(1138) + adder_tree(0)(1139); --27 bits 
            adder_tree(1)(570) <= adder_tree(0)(1140) + adder_tree(0)(1141); --27 bits 
            adder_tree(1)(571) <= adder_tree(0)(1142) + adder_tree(0)(1143); --27 bits 
            adder_tree(1)(572) <= adder_tree(0)(1144) + adder_tree(0)(1145); --27 bits 
            adder_tree(1)(573) <= adder_tree(0)(1146) + adder_tree(0)(1147); --27 bits 
            adder_tree(1)(574) <= adder_tree(0)(1148) + adder_tree(0)(1149); --27 bits 
            adder_tree(1)(575) <= adder_tree(0)(1150) + adder_tree(0)(1151); --27 bits 
            adder_tree(1)(576) <= adder_tree(0)(1152) + adder_tree(0)(1153); --27 bits 
            adder_tree(1)(577) <= adder_tree(0)(1154) + adder_tree(0)(1155); --27 bits 
            adder_tree(1)(578) <= adder_tree(0)(1156) + adder_tree(0)(1157); --27 bits 
            adder_tree(1)(579) <= adder_tree(0)(1158) + adder_tree(0)(1159); --27 bits 
            adder_tree(1)(580) <= adder_tree(0)(1160) + adder_tree(0)(1161); --27 bits 
            adder_tree(1)(581) <= adder_tree(0)(1162) + adder_tree(0)(1163); --27 bits 
            adder_tree(1)(582) <= adder_tree(0)(1164) + adder_tree(0)(1165); --27 bits 
            adder_tree(1)(583) <= adder_tree(0)(1166) + adder_tree(0)(1167); --27 bits 
            adder_tree(1)(584) <= adder_tree(0)(1168) + adder_tree(0)(1169); --27 bits 
            adder_tree(1)(585) <= adder_tree(0)(1170) + adder_tree(0)(1171); --27 bits 
            adder_tree(1)(586) <= adder_tree(0)(1172) + adder_tree(0)(1173); --27 bits 
            adder_tree(1)(587) <= adder_tree(0)(1174) + adder_tree(0)(1175); --27 bits 
            adder_tree(1)(588) <= adder_tree(0)(1176) + adder_tree(0)(1177); --27 bits 
            adder_tree(1)(589) <= adder_tree(0)(1178) + adder_tree(0)(1179); --27 bits 
            adder_tree(1)(590) <= adder_tree(0)(1180) + adder_tree(0)(1181); --27 bits 
            adder_tree(1)(591) <= adder_tree(0)(1182) + adder_tree(0)(1183); --27 bits 
            adder_tree(1)(592) <= adder_tree(0)(1184) + adder_tree(0)(1185); --27 bits 
            adder_tree(1)(593) <= adder_tree(0)(1186) + adder_tree(0)(1187); --27 bits 
            adder_tree(1)(594) <= adder_tree(0)(1188) + adder_tree(0)(1189); --27 bits 
            adder_tree(1)(595) <= adder_tree(0)(1190) + adder_tree(0)(1191); --27 bits 
            adder_tree(1)(596) <= adder_tree(0)(1192) + adder_tree(0)(1193); --27 bits 
            adder_tree(1)(597) <= adder_tree(0)(1194) + adder_tree(0)(1195); --27 bits 
            adder_tree(1)(598) <= adder_tree(0)(1196) + adder_tree(0)(1197); --27 bits 
            adder_tree(1)(599) <= adder_tree(0)(1198) + adder_tree(0)(1199); --27 bits 
            adder_tree(1)(600) <= adder_tree(0)(1200) + adder_tree(0)(1201); --27 bits 
            adder_tree(1)(601) <= adder_tree(0)(1202) + adder_tree(0)(1203); --27 bits 
            adder_tree(1)(602) <= adder_tree(0)(1204) + adder_tree(0)(1205); --27 bits 
            adder_tree(1)(603) <= adder_tree(0)(1206) + adder_tree(0)(1207); --27 bits 
            adder_tree(1)(604) <= adder_tree(0)(1208) + adder_tree(0)(1209); --27 bits 
            adder_tree(1)(605) <= adder_tree(0)(1210) + adder_tree(0)(1211); --27 bits 
            adder_tree(1)(606) <= adder_tree(0)(1212) + adder_tree(0)(1213); --27 bits 
            adder_tree(1)(607) <= adder_tree(0)(1214) + adder_tree(0)(1215); --27 bits 
            adder_tree(1)(608) <= adder_tree(0)(1216) + adder_tree(0)(1217); --27 bits 
            adder_tree(1)(609) <= adder_tree(0)(1218) + adder_tree(0)(1219); --27 bits 
            adder_tree(1)(610) <= adder_tree(0)(1220) + adder_tree(0)(1221); --27 bits 
            adder_tree(1)(611) <= adder_tree(0)(1222) + adder_tree(0)(1223); --27 bits 
            adder_tree(1)(612) <= adder_tree(0)(1224) + adder_tree(0)(1225); --27 bits 
            adder_tree(1)(613) <= adder_tree(0)(1226) + adder_tree(0)(1227); --27 bits 
            adder_tree(1)(614) <= adder_tree(0)(1228) + adder_tree(0)(1229); --27 bits 
            adder_tree(1)(615) <= adder_tree(0)(1230) + adder_tree(0)(1231); --27 bits 
            adder_tree(1)(616) <= adder_tree(0)(1232) + adder_tree(0)(1233); --27 bits 
            adder_tree(1)(617) <= adder_tree(0)(1234) + adder_tree(0)(1235); --27 bits 
            adder_tree(1)(618) <= adder_tree(0)(1236) + adder_tree(0)(1237); --27 bits 
            adder_tree(1)(619) <= adder_tree(0)(1238) + adder_tree(0)(1239); --27 bits 
            adder_tree(1)(620) <= adder_tree(0)(1240) + adder_tree(0)(1241); --27 bits 
            adder_tree(1)(621) <= adder_tree(0)(1242) + adder_tree(0)(1243); --27 bits 
            adder_tree(1)(622) <= adder_tree(0)(1244) + adder_tree(0)(1245); --27 bits 
            adder_tree(1)(623) <= adder_tree(0)(1246) + adder_tree(0)(1247); --27 bits 
            adder_tree(1)(624) <= adder_tree(0)(1248) + adder_tree(0)(1249); --27 bits 
            adder_tree(1)(625) <= adder_tree(0)(1250) + adder_tree(0)(1251); --27 bits 
            adder_tree(1)(626) <= adder_tree(0)(1252) + adder_tree(0)(1253); --27 bits 
            adder_tree(1)(627) <= adder_tree(0)(1254) + adder_tree(0)(1255); --27 bits 
            adder_tree(1)(628) <= adder_tree(0)(1256) + adder_tree(0)(1257); --27 bits 
            adder_tree(1)(629) <= adder_tree(0)(1258) + adder_tree(0)(1259); --27 bits 
            adder_tree(1)(630) <= adder_tree(0)(1260) + adder_tree(0)(1261); --27 bits 
            adder_tree(1)(631) <= adder_tree(0)(1262) + adder_tree(0)(1263); --27 bits 
            adder_tree(1)(632) <= adder_tree(0)(1264) + adder_tree(0)(1265); --27 bits 
            adder_tree(1)(633) <= adder_tree(0)(1266) + adder_tree(0)(1267); --27 bits 
            adder_tree(1)(634) <= adder_tree(0)(1268) + adder_tree(0)(1269); --27 bits 
            adder_tree(1)(635) <= adder_tree(0)(1270) + adder_tree(0)(1271); --27 bits 
            adder_tree(1)(636) <= adder_tree(0)(1272) + adder_tree(0)(1273); --27 bits 
            adder_tree(1)(637) <= adder_tree(0)(1274) + adder_tree(0)(1275); --27 bits 
            adder_tree(1)(638) <= adder_tree(0)(1276) + adder_tree(0)(1277); --27 bits 
            adder_tree(1)(639) <= adder_tree(0)(1278) + adder_tree(0)(1279); --27 bits 
            adder_tree(1)(640) <= adder_tree(0)(1280) + adder_tree(0)(1281); --27 bits 
            adder_tree(1)(641) <= adder_tree(0)(1282) + adder_tree(0)(1283); --27 bits 
            adder_tree(1)(642) <= adder_tree(0)(1284) + adder_tree(0)(1285); --27 bits 
            adder_tree(1)(643) <= adder_tree(0)(1286) + adder_tree(0)(1287); --27 bits 
            adder_tree(1)(644) <= adder_tree(0)(1288) + adder_tree(0)(1289); --27 bits 
            adder_tree(1)(645) <= adder_tree(0)(1290) + adder_tree(0)(1291); --27 bits 
            adder_tree(1)(646) <= adder_tree(0)(1292) + adder_tree(0)(1293); --27 bits 
            adder_tree(1)(647) <= adder_tree(0)(1294) + adder_tree(0)(1295); --27 bits 
            adder_tree(1)(648) <= adder_tree(0)(1296) + adder_tree(0)(1297); --27 bits 
            adder_tree(1)(649) <= adder_tree(0)(1298) + adder_tree(0)(1299); --27 bits 
            adder_tree(1)(650) <= adder_tree(0)(1300) + adder_tree(0)(1301); --27 bits 
            adder_tree(1)(651) <= adder_tree(0)(1302) + adder_tree(0)(1303); --27 bits 
            adder_tree(1)(652) <= adder_tree(0)(1304) + adder_tree(0)(1305); --27 bits 
            adder_tree(1)(653) <= adder_tree(0)(1306) + adder_tree(0)(1307); --27 bits 
            adder_tree(1)(654) <= adder_tree(0)(1308) + adder_tree(0)(1309); --27 bits 
            adder_tree(1)(655) <= adder_tree(0)(1310) + adder_tree(0)(1311); --27 bits 
            adder_tree(1)(656) <= adder_tree(0)(1312) + adder_tree(0)(1313); --27 bits 
            adder_tree(1)(657) <= adder_tree(0)(1314) + adder_tree(0)(1315); --27 bits 
            adder_tree(1)(658) <= adder_tree(0)(1316) + adder_tree(0)(1317); --27 bits 
            adder_tree(1)(659) <= adder_tree(0)(1318) + adder_tree(0)(1319); --27 bits 
            adder_tree(1)(660) <= adder_tree(0)(1320) + adder_tree(0)(1321); --27 bits 
            adder_tree(1)(661) <= adder_tree(0)(1322) + adder_tree(0)(1323); --27 bits 
            adder_tree(1)(662) <= adder_tree(0)(1324) + adder_tree(0)(1325); --27 bits 
            adder_tree(1)(663) <= adder_tree(0)(1326) + adder_tree(0)(1327); --27 bits 
            adder_tree(1)(664) <= adder_tree(0)(1328) + adder_tree(0)(1329); --27 bits 
            adder_tree(1)(665) <= adder_tree(0)(1330) + adder_tree(0)(1331); --27 bits 
            adder_tree(1)(666) <= adder_tree(0)(1332) + adder_tree(0)(1333); --27 bits 
            adder_tree(1)(667) <= adder_tree(0)(1334) + adder_tree(0)(1335); --27 bits 
            adder_tree(1)(668) <= adder_tree(0)(1336) + adder_tree(0)(1337); --27 bits 
            adder_tree(1)(669) <= adder_tree(0)(1338) + adder_tree(0)(1339); --27 bits 
            adder_tree(1)(670) <= adder_tree(0)(1340) + adder_tree(0)(1341); --27 bits 
            adder_tree(1)(671) <= adder_tree(0)(1342) + adder_tree(0)(1343); --27 bits 
            adder_tree(1)(672) <= adder_tree(0)(1344) + adder_tree(0)(1345); --27 bits 
            adder_tree(1)(673) <= adder_tree(0)(1346) + adder_tree(0)(1347); --27 bits 
            adder_tree(1)(674) <= adder_tree(0)(1348) + adder_tree(0)(1349); --27 bits 
            adder_tree(1)(675) <= adder_tree(0)(1350) + adder_tree(0)(1351); --27 bits 
            adder_tree(1)(676) <= adder_tree(0)(1352) + adder_tree(0)(1353); --27 bits 
            adder_tree(1)(677) <= adder_tree(0)(1354) + adder_tree(0)(1355); --27 bits 
            adder_tree(1)(678) <= adder_tree(0)(1356) + adder_tree(0)(1357); --27 bits 
            adder_tree(1)(679) <= adder_tree(0)(1358) + adder_tree(0)(1359); --27 bits 
            adder_tree(1)(680) <= adder_tree(0)(1360) + adder_tree(0)(1361); --27 bits 
            adder_tree(1)(681) <= adder_tree(0)(1362) + adder_tree(0)(1363); --27 bits 
            adder_tree(1)(682) <= adder_tree(0)(1364) + adder_tree(0)(1365); --27 bits 
            adder_tree(1)(683) <= adder_tree(0)(1366) + adder_tree(0)(1367); --27 bits 
            adder_tree(1)(684) <= adder_tree(0)(1368) + adder_tree(0)(1369); --27 bits 
            adder_tree(1)(685) <= adder_tree(0)(1370) + adder_tree(0)(1371); --27 bits 
            adder_tree(1)(686) <= adder_tree(0)(1372) + adder_tree(0)(1373); --27 bits 
            adder_tree(1)(687) <= adder_tree(0)(1374) + adder_tree(0)(1375); --27 bits 
            adder_tree(1)(688) <= adder_tree(0)(1376) + adder_tree(0)(1377); --27 bits 
            adder_tree(1)(689) <= adder_tree(0)(1378) + adder_tree(0)(1379); --27 bits 
            adder_tree(1)(690) <= adder_tree(0)(1380) + adder_tree(0)(1381); --27 bits 
            adder_tree(1)(691) <= adder_tree(0)(1382) + adder_tree(0)(1383); --27 bits 
            adder_tree(1)(692) <= adder_tree(0)(1384) + adder_tree(0)(1385); --27 bits 
            adder_tree(1)(693) <= adder_tree(0)(1386) + adder_tree(0)(1387); --27 bits 
            adder_tree(1)(694) <= adder_tree(0)(1388) + adder_tree(0)(1389); --27 bits 
            adder_tree(1)(695) <= adder_tree(0)(1390) + adder_tree(0)(1391); --27 bits 
            adder_tree(1)(696) <= adder_tree(0)(1392) + adder_tree(0)(1393); --27 bits 
            adder_tree(1)(697) <= adder_tree(0)(1394) + adder_tree(0)(1395); --27 bits 
            adder_tree(1)(698) <= adder_tree(0)(1396) + adder_tree(0)(1397); --27 bits 
            adder_tree(1)(699) <= adder_tree(0)(1398) + adder_tree(0)(1399); --27 bits 
            adder_tree(1)(700) <= adder_tree(0)(1400) + adder_tree(0)(1401); --27 bits 
            adder_tree(1)(701) <= adder_tree(0)(1402) + adder_tree(0)(1403); --27 bits 
            adder_tree(1)(702) <= adder_tree(0)(1404) + adder_tree(0)(1405); --27 bits 
            adder_tree(1)(703) <= adder_tree(0)(1406) + adder_tree(0)(1407); --27 bits 
            adder_tree(1)(704) <= adder_tree(0)(1408) + adder_tree(0)(1409); --27 bits 
            adder_tree(1)(705) <= adder_tree(0)(1410) + adder_tree(0)(1411); --27 bits 
            adder_tree(1)(706) <= adder_tree(0)(1412) + adder_tree(0)(1413); --27 bits 
            adder_tree(1)(707) <= adder_tree(0)(1414) + adder_tree(0)(1415); --27 bits 
            adder_tree(1)(708) <= adder_tree(0)(1416) + adder_tree(0)(1417); --27 bits 
            adder_tree(1)(709) <= adder_tree(0)(1418) + adder_tree(0)(1419); --27 bits 
            adder_tree(1)(710) <= adder_tree(0)(1420) + adder_tree(0)(1421); --27 bits 
            adder_tree(1)(711) <= adder_tree(0)(1422) + adder_tree(0)(1423); --27 bits 
            adder_tree(1)(712) <= adder_tree(0)(1424) + adder_tree(0)(1425); --27 bits 
            adder_tree(1)(713) <= adder_tree(0)(1426) + adder_tree(0)(1427); --27 bits 
            adder_tree(1)(714) <= adder_tree(0)(1428) + adder_tree(0)(1429); --27 bits 
            adder_tree(1)(715) <= adder_tree(0)(1430) + adder_tree(0)(1431); --27 bits 
            adder_tree(1)(716) <= adder_tree(0)(1432) + adder_tree(0)(1433); --27 bits 
            adder_tree(1)(717) <= adder_tree(0)(1434) + adder_tree(0)(1435); --27 bits 
            adder_tree(1)(718) <= adder_tree(0)(1436) + adder_tree(0)(1437); --27 bits 
            adder_tree(1)(719) <= adder_tree(0)(1438) + adder_tree(0)(1439); --27 bits 
            adder_tree(1)(720) <= adder_tree(0)(1440) + adder_tree(0)(1441); --27 bits 
            adder_tree(1)(721) <= adder_tree(0)(1442) + adder_tree(0)(1443); --27 bits 
            adder_tree(1)(722) <= adder_tree(0)(1444) + adder_tree(0)(1445); --27 bits 
            adder_tree(1)(723) <= adder_tree(0)(1446) + adder_tree(0)(1447); --27 bits 
            adder_tree(1)(724) <= adder_tree(0)(1448) + adder_tree(0)(1449); --27 bits 
            adder_tree(1)(725) <= adder_tree(0)(1450) + adder_tree(0)(1451); --27 bits 
            adder_tree(1)(726) <= adder_tree(0)(1452) + adder_tree(0)(1453); --27 bits 
            adder_tree(1)(727) <= adder_tree(0)(1454) + adder_tree(0)(1455); --27 bits 
            adder_tree(1)(728) <= adder_tree(0)(1456) + adder_tree(0)(1457); --27 bits 
            adder_tree(1)(729) <= adder_tree(0)(1458) + adder_tree(0)(1459); --27 bits 
            adder_tree(1)(730) <= adder_tree(0)(1460) + adder_tree(0)(1461); --27 bits 
            adder_tree(1)(731) <= adder_tree(0)(1462) + adder_tree(0)(1463); --27 bits 
            adder_tree(1)(732) <= adder_tree(0)(1464) + adder_tree(0)(1465); --27 bits 
            adder_tree(1)(733) <= adder_tree(0)(1466) + adder_tree(0)(1467); --27 bits 
            adder_tree(1)(734) <= adder_tree(0)(1468) + adder_tree(0)(1469); --27 bits 
            adder_tree(1)(735) <= adder_tree(0)(1470) + adder_tree(0)(1471); --27 bits 
            adder_tree(1)(736) <= adder_tree(0)(1472) + adder_tree(0)(1473); --27 bits 
            adder_tree(1)(737) <= adder_tree(0)(1474) + adder_tree(0)(1475); --27 bits 
            adder_tree(1)(738) <= adder_tree(0)(1476) + adder_tree(0)(1477); --27 bits 
            adder_tree(1)(739) <= adder_tree(0)(1478) + adder_tree(0)(1479); --27 bits 
            adder_tree(1)(740) <= adder_tree(0)(1480) + adder_tree(0)(1481); --27 bits 
            adder_tree(1)(741) <= adder_tree(0)(1482) + adder_tree(0)(1483); --27 bits 
            adder_tree(1)(742) <= adder_tree(0)(1484) + adder_tree(0)(1485); --27 bits 
            adder_tree(1)(743) <= adder_tree(0)(1486) + adder_tree(0)(1487); --27 bits 
            adder_tree(1)(744) <= adder_tree(0)(1488) + adder_tree(0)(1489); --27 bits 
            adder_tree(1)(745) <= adder_tree(0)(1490) + adder_tree(0)(1491); --27 bits 
            adder_tree(1)(746) <= adder_tree(0)(1492) + adder_tree(0)(1493); --27 bits 
            adder_tree(1)(747) <= adder_tree(0)(1494) + adder_tree(0)(1495); --27 bits 
            adder_tree(1)(748) <= adder_tree(0)(1496) + adder_tree(0)(1497); --27 bits 
            adder_tree(1)(749) <= adder_tree(0)(1498) + adder_tree(0)(1499); --27 bits 
            adder_tree(1)(750) <= adder_tree(0)(1500) + adder_tree(0)(1501); --27 bits 
            adder_tree(1)(751) <= adder_tree(0)(1502) + adder_tree(0)(1503); --27 bits 
            adder_tree(1)(752) <= adder_tree(0)(1504) + adder_tree(0)(1505); --27 bits 
            adder_tree(1)(753) <= adder_tree(0)(1506) + adder_tree(0)(1507); --27 bits 
            adder_tree(1)(754) <= adder_tree(0)(1508) + adder_tree(0)(1509); --27 bits 
            adder_tree(1)(755) <= adder_tree(0)(1510) + adder_tree(0)(1511); --27 bits 
            adder_tree(1)(756) <= adder_tree(0)(1512) + adder_tree(0)(1513); --27 bits 
            adder_tree(1)(757) <= adder_tree(0)(1514) + adder_tree(0)(1515); --27 bits 
            adder_tree(1)(758) <= adder_tree(0)(1516) + adder_tree(0)(1517); --27 bits 
            adder_tree(1)(759) <= adder_tree(0)(1518) + adder_tree(0)(1519); --27 bits 
            adder_tree(1)(760) <= adder_tree(0)(1520) + adder_tree(0)(1521); --27 bits 
            adder_tree(1)(761) <= adder_tree(0)(1522) + adder_tree(0)(1523); --27 bits 
            adder_tree(1)(762) <= adder_tree(0)(1524) + adder_tree(0)(1525); --27 bits 
            adder_tree(1)(763) <= adder_tree(0)(1526) + adder_tree(0)(1527); --27 bits 
            adder_tree(1)(764) <= adder_tree(0)(1528) + adder_tree(0)(1529); --27 bits 
            adder_tree(1)(765) <= adder_tree(0)(1530) + adder_tree(0)(1531); --27 bits 
            adder_tree(1)(766) <= adder_tree(0)(1532) + adder_tree(0)(1533); --27 bits 
            adder_tree(1)(767) <= adder_tree(0)(1534) + adder_tree(0)(1535); --27 bits 
            adder_tree(1)(768) <= adder_tree(0)(1536) + adder_tree(0)(1537); --27 bits 
            adder_tree(1)(769) <= adder_tree(0)(1538) + adder_tree(0)(1539); --27 bits 
            adder_tree(1)(770) <= adder_tree(0)(1540) + adder_tree(0)(1541); --27 bits 
            adder_tree(1)(771) <= adder_tree(0)(1542) + adder_tree(0)(1543); --27 bits 
            adder_tree(1)(772) <= adder_tree(0)(1544) + adder_tree(0)(1545); --27 bits 
            adder_tree(1)(773) <= adder_tree(0)(1546) + adder_tree(0)(1547); --27 bits 
            adder_tree(1)(774) <= adder_tree(0)(1548) + adder_tree(0)(1549); --27 bits 
            adder_tree(1)(775) <= adder_tree(0)(1550) + adder_tree(0)(1551); --27 bits 
            adder_tree(1)(776) <= adder_tree(0)(1552) + adder_tree(0)(1553); --27 bits 
            adder_tree(1)(777) <= adder_tree(0)(1554) + adder_tree(0)(1555); --27 bits 
            adder_tree(1)(778) <= adder_tree(0)(1556) + adder_tree(0)(1557); --27 bits 
            adder_tree(1)(779) <= adder_tree(0)(1558) + adder_tree(0)(1559); --27 bits 
            adder_tree(1)(780) <= adder_tree(0)(1560) + adder_tree(0)(1561); --27 bits 
            adder_tree(1)(781) <= adder_tree(0)(1562) + adder_tree(0)(1563); --27 bits 
            adder_tree(1)(782) <= adder_tree(0)(1564) + adder_tree(0)(1565); --27 bits 
            adder_tree(1)(783) <= adder_tree(0)(1566) + adder_tree(0)(1567); --27 bits 
            adder_tree(1)(784) <= adder_tree(0)(1568) + adder_tree(0)(1569); --27 bits 
            adder_tree(1)(785) <= adder_tree(0)(1570) + adder_tree(0)(1571); --27 bits 
            adder_tree(1)(786) <= adder_tree(0)(1572) + adder_tree(0)(1573); --27 bits 
            adder_tree(1)(787) <= adder_tree(0)(1574) + adder_tree(0)(1575); --27 bits 
            adder_tree(1)(788) <= adder_tree(0)(1576) + adder_tree(0)(1577); --27 bits 
            adder_tree(1)(789) <= adder_tree(0)(1578) + adder_tree(0)(1579); --27 bits 
            adder_tree(1)(790) <= adder_tree(0)(1580) + adder_tree(0)(1581); --27 bits 
            adder_tree(1)(791) <= adder_tree(0)(1582) + adder_tree(0)(1583); --27 bits 
            adder_tree(1)(792) <= adder_tree(0)(1584) + adder_tree(0)(1585); --27 bits 
            adder_tree(1)(793) <= adder_tree(0)(1586) + adder_tree(0)(1587); --27 bits 
            adder_tree(1)(794) <= adder_tree(0)(1588) + adder_tree(0)(1589); --27 bits 
            adder_tree(1)(795) <= adder_tree(0)(1590) + adder_tree(0)(1591); --27 bits 
            adder_tree(1)(796) <= adder_tree(0)(1592) + adder_tree(0)(1593); --27 bits 
            adder_tree(1)(797) <= adder_tree(0)(1594) + adder_tree(0)(1595); --27 bits 
            adder_tree(1)(798) <= adder_tree(0)(1596) + adder_tree(0)(1597); --27 bits 
            adder_tree(1)(799) <= adder_tree(0)(1598) + adder_tree(0)(1599); --27 bits 
            adder_tree(1)(800) <= adder_tree(0)(1600) + adder_tree(0)(1601); --27 bits 
            adder_tree(1)(801) <= adder_tree(0)(1602) + adder_tree(0)(1603); --27 bits 
            adder_tree(1)(802) <= adder_tree(0)(1604) + adder_tree(0)(1605); --27 bits 
            adder_tree(1)(803) <= adder_tree(0)(1606) + adder_tree(0)(1607); --27 bits 
            adder_tree(1)(804) <= adder_tree(0)(1608) + adder_tree(0)(1609); --27 bits 
            adder_tree(1)(805) <= adder_tree(0)(1610) + adder_tree(0)(1611); --27 bits 
            adder_tree(1)(806) <= adder_tree(0)(1612) + adder_tree(0)(1613); --27 bits 
            adder_tree(1)(807) <= adder_tree(0)(1614) + adder_tree(0)(1615); --27 bits 
            adder_tree(1)(808) <= adder_tree(0)(1616) + adder_tree(0)(1617); --27 bits 
            adder_tree(1)(809) <= adder_tree(0)(1618) + adder_tree(0)(1619); --27 bits 
            adder_tree(1)(810) <= adder_tree(0)(1620) + adder_tree(0)(1621); --27 bits 
            adder_tree(1)(811) <= adder_tree(0)(1622) + adder_tree(0)(1623); --27 bits 
            adder_tree(1)(812) <= adder_tree(0)(1624) + adder_tree(0)(1625); --27 bits 
            adder_tree(1)(813) <= adder_tree(0)(1626) + adder_tree(0)(1627); --27 bits 
            adder_tree(1)(814) <= adder_tree(0)(1628) + adder_tree(0)(1629); --27 bits 
            adder_tree(1)(815) <= adder_tree(0)(1630) + adder_tree(0)(1631); --27 bits 
            adder_tree(1)(816) <= adder_tree(0)(1632) + adder_tree(0)(1633); --27 bits 
            adder_tree(1)(817) <= adder_tree(0)(1634) + adder_tree(0)(1635); --27 bits 
            adder_tree(1)(818) <= adder_tree(0)(1636) + adder_tree(0)(1637); --27 bits 
            adder_tree(1)(819) <= adder_tree(0)(1638) + adder_tree(0)(1639); --27 bits 
            adder_tree(1)(820) <= adder_tree(0)(1640) + adder_tree(0)(1641); --27 bits 
            adder_tree(1)(821) <= adder_tree(0)(1642) + adder_tree(0)(1643); --27 bits 
            adder_tree(1)(822) <= adder_tree(0)(1644) + adder_tree(0)(1645); --27 bits 
            adder_tree(1)(823) <= adder_tree(0)(1646) + adder_tree(0)(1647); --27 bits 
            adder_tree(1)(824) <= adder_tree(0)(1648) + adder_tree(0)(1649); --27 bits 
            adder_tree(1)(825) <= adder_tree(0)(1650) + adder_tree(0)(1651); --27 bits 
            adder_tree(1)(826) <= adder_tree(0)(1652) + adder_tree(0)(1653); --27 bits 
            adder_tree(1)(827) <= adder_tree(0)(1654) + adder_tree(0)(1655); --27 bits 
            adder_tree(1)(828) <= adder_tree(0)(1656) + adder_tree(0)(1657); --27 bits 
            adder_tree(1)(829) <= adder_tree(0)(1658) + adder_tree(0)(1659); --27 bits 
            adder_tree(1)(830) <= adder_tree(0)(1660) + adder_tree(0)(1661); --27 bits 
            adder_tree(1)(831) <= adder_tree(0)(1662) + adder_tree(0)(1663); --27 bits 
            adder_tree(1)(832) <= adder_tree(0)(1664) + adder_tree(0)(1665); --27 bits 
            adder_tree(1)(833) <= adder_tree(0)(1666) + adder_tree(0)(1667); --27 bits 
            adder_tree(1)(834) <= adder_tree(0)(1668) + adder_tree(0)(1669); --27 bits 
            adder_tree(1)(835) <= adder_tree(0)(1670) + adder_tree(0)(1671); --27 bits 
            adder_tree(1)(836) <= adder_tree(0)(1672) + adder_tree(0)(1673); --27 bits 
            adder_tree(1)(837) <= adder_tree(0)(1674) + adder_tree(0)(1675); --27 bits 
            adder_tree(1)(838) <= adder_tree(0)(1676) + adder_tree(0)(1677); --27 bits 
            adder_tree(1)(839) <= adder_tree(0)(1678) + adder_tree(0)(1679); --27 bits 
            adder_tree(1)(840) <= adder_tree(0)(1680) + adder_tree(0)(1681); --27 bits 
            adder_tree(1)(841) <= adder_tree(0)(1682) + adder_tree(0)(1683); --27 bits 
            adder_tree(1)(842) <= adder_tree(0)(1684) + adder_tree(0)(1685); --27 bits 
            adder_tree(1)(843) <= adder_tree(0)(1686) + adder_tree(0)(1687); --27 bits 
            adder_tree(1)(844) <= adder_tree(0)(1688) + adder_tree(0)(1689); --27 bits 
            adder_tree(1)(845) <= adder_tree(0)(1690) + adder_tree(0)(1691); --27 bits 
            adder_tree(1)(846) <= adder_tree(0)(1692) + adder_tree(0)(1693); --27 bits 
            adder_tree(1)(847) <= adder_tree(0)(1694) + adder_tree(0)(1695); --27 bits 
            adder_tree(1)(848) <= adder_tree(0)(1696) + adder_tree(0)(1697); --27 bits 
            adder_tree(1)(849) <= adder_tree(0)(1698) + adder_tree(0)(1699); --27 bits 
            adder_tree(1)(850) <= adder_tree(0)(1700) + adder_tree(0)(1701); --27 bits 
            adder_tree(1)(851) <= adder_tree(0)(1702) + adder_tree(0)(1703); --27 bits 
            adder_tree(1)(852) <= adder_tree(0)(1704) + adder_tree(0)(1705); --27 bits 
            adder_tree(1)(853) <= adder_tree(0)(1706) + adder_tree(0)(1707); --27 bits 
            adder_tree(1)(854) <= adder_tree(0)(1708) + adder_tree(0)(1709); --27 bits 
            adder_tree(1)(855) <= adder_tree(0)(1710) + adder_tree(0)(1711); --27 bits 
            adder_tree(1)(856) <= adder_tree(0)(1712) + adder_tree(0)(1713); --27 bits 
            adder_tree(1)(857) <= adder_tree(0)(1714) + adder_tree(0)(1715); --27 bits 
            adder_tree(1)(858) <= adder_tree(0)(1716) + adder_tree(0)(1717); --27 bits 
            adder_tree(1)(859) <= adder_tree(0)(1718) + adder_tree(0)(1719); --27 bits 
            adder_tree(1)(860) <= adder_tree(0)(1720) + adder_tree(0)(1721); --27 bits 
            adder_tree(1)(861) <= adder_tree(0)(1722) + adder_tree(0)(1723); --27 bits 
            adder_tree(1)(862) <= adder_tree(0)(1724) + adder_tree(0)(1725); --27 bits 
            adder_tree(1)(863) <= adder_tree(0)(1726) + adder_tree(0)(1727); --27 bits 
            adder_tree(1)(864) <= adder_tree(0)(1728) + adder_tree(0)(1729); --27 bits 
            adder_tree(1)(865) <= adder_tree(0)(1730) + adder_tree(0)(1731); --27 bits 
            adder_tree(1)(866) <= adder_tree(0)(1732) + adder_tree(0)(1733); --27 bits 
            adder_tree(1)(867) <= adder_tree(0)(1734) + adder_tree(0)(1735); --27 bits 
            adder_tree(1)(868) <= adder_tree(0)(1736) + adder_tree(0)(1737); --27 bits 
            adder_tree(1)(869) <= adder_tree(0)(1738) + adder_tree(0)(1739); --27 bits 
            adder_tree(1)(870) <= adder_tree(0)(1740) + adder_tree(0)(1741); --27 bits 
            adder_tree(1)(871) <= adder_tree(0)(1742) + adder_tree(0)(1743); --27 bits 
            adder_tree(1)(872) <= adder_tree(0)(1744) + adder_tree(0)(1745); --27 bits 
            adder_tree(1)(873) <= adder_tree(0)(1746) + adder_tree(0)(1747); --27 bits 
            adder_tree(1)(874) <= adder_tree(0)(1748) + adder_tree(0)(1749); --27 bits 
            adder_tree(1)(875) <= adder_tree(0)(1750) + adder_tree(0)(1751); --27 bits 
            adder_tree(1)(876) <= adder_tree(0)(1752) + adder_tree(0)(1753); --27 bits 
            adder_tree(1)(877) <= adder_tree(0)(1754) + adder_tree(0)(1755); --27 bits 
            adder_tree(1)(878) <= adder_tree(0)(1756) + adder_tree(0)(1757); --27 bits 
            adder_tree(1)(879) <= adder_tree(0)(1758) + adder_tree(0)(1759); --27 bits 
            adder_tree(1)(880) <= adder_tree(0)(1760) + adder_tree(0)(1761); --27 bits 
            adder_tree(1)(881) <= adder_tree(0)(1762) + adder_tree(0)(1763); --27 bits 
            adder_tree(1)(882) <= adder_tree(0)(1764) + adder_tree(0)(1765); --27 bits 
            adder_tree(1)(883) <= adder_tree(0)(1766) + adder_tree(0)(1767); --27 bits 
            adder_tree(1)(884) <= adder_tree(0)(1768) + adder_tree(0)(1769); --27 bits 
            adder_tree(1)(885) <= adder_tree(0)(1770) + adder_tree(0)(1771); --27 bits 
            adder_tree(1)(886) <= adder_tree(0)(1772) + adder_tree(0)(1773); --27 bits 
            adder_tree(1)(887) <= adder_tree(0)(1774) + adder_tree(0)(1775); --27 bits 
            adder_tree(1)(888) <= adder_tree(0)(1776) + adder_tree(0)(1777); --27 bits 
            adder_tree(1)(889) <= adder_tree(0)(1778) + adder_tree(0)(1779); --27 bits 
            adder_tree(1)(890) <= adder_tree(0)(1780) + adder_tree(0)(1781); --27 bits 
            adder_tree(1)(891) <= adder_tree(0)(1782) + adder_tree(0)(1783); --27 bits 
            adder_tree(1)(892) <= adder_tree(0)(1784) + adder_tree(0)(1785); --27 bits 
            adder_tree(1)(893) <= adder_tree(0)(1786) + adder_tree(0)(1787); --27 bits 
            adder_tree(1)(894) <= adder_tree(0)(1788) + adder_tree(0)(1789); --27 bits 
            adder_tree(1)(895) <= adder_tree(0)(1790) + adder_tree(0)(1791); --27 bits 
            adder_tree(1)(896) <= adder_tree(0)(1792) + adder_tree(0)(1793); --27 bits 
            adder_tree(1)(897) <= adder_tree(0)(1794) + adder_tree(0)(1795); --27 bits 
            adder_tree(1)(898) <= adder_tree(0)(1796) + adder_tree(0)(1797); --27 bits 
            adder_tree(1)(899) <= adder_tree(0)(1798) + adder_tree(0)(1799); --27 bits 
            adder_tree(1)(900) <= adder_tree(0)(1800) + adder_tree(0)(1801); --27 bits 
            adder_tree(1)(901) <= adder_tree(0)(1802) + adder_tree(0)(1803); --27 bits 
            adder_tree(1)(902) <= adder_tree(0)(1804) + adder_tree(0)(1805); --27 bits 
            adder_tree(1)(903) <= adder_tree(0)(1806) + adder_tree(0)(1807); --27 bits 
            adder_tree(1)(904) <= adder_tree(0)(1808) + adder_tree(0)(1809); --27 bits 
            adder_tree(1)(905) <= adder_tree(0)(1810) + adder_tree(0)(1811); --27 bits 
            adder_tree(1)(906) <= adder_tree(0)(1812) + adder_tree(0)(1813); --27 bits 
            adder_tree(1)(907) <= adder_tree(0)(1814) + adder_tree(0)(1815); --27 bits 
            adder_tree(1)(908) <= adder_tree(0)(1816) + adder_tree(0)(1817); --27 bits 
            adder_tree(1)(909) <= adder_tree(0)(1818) + adder_tree(0)(1819); --27 bits 
            adder_tree(1)(910) <= adder_tree(0)(1820) + adder_tree(0)(1821); --27 bits 
            adder_tree(1)(911) <= adder_tree(0)(1822) + adder_tree(0)(1823); --27 bits 
            adder_tree(1)(912) <= adder_tree(0)(1824) + adder_tree(0)(1825); --27 bits 
            adder_tree(1)(913) <= adder_tree(0)(1826) + adder_tree(0)(1827); --27 bits 
            adder_tree(1)(914) <= adder_tree(0)(1828) + adder_tree(0)(1829); --27 bits 
            adder_tree(1)(915) <= adder_tree(0)(1830) + adder_tree(0)(1831); --27 bits 
            adder_tree(1)(916) <= adder_tree(0)(1832) + adder_tree(0)(1833); --27 bits 
            adder_tree(1)(917) <= adder_tree(0)(1834) + adder_tree(0)(1835); --27 bits 
            adder_tree(1)(918) <= adder_tree(0)(1836) + adder_tree(0)(1837); --27 bits 
            adder_tree(1)(919) <= adder_tree(0)(1838) + adder_tree(0)(1839); --27 bits 
            adder_tree(1)(920) <= adder_tree(0)(1840) + adder_tree(0)(1841); --27 bits 
            adder_tree(1)(921) <= adder_tree(0)(1842) + adder_tree(0)(1843); --27 bits 
            adder_tree(1)(922) <= adder_tree(0)(1844) + adder_tree(0)(1845); --27 bits 
            adder_tree(1)(923) <= adder_tree(0)(1846) + adder_tree(0)(1847); --27 bits 
            adder_tree(1)(924) <= adder_tree(0)(1848) + adder_tree(0)(1849); --27 bits 
            adder_tree(1)(925) <= adder_tree(0)(1850) + adder_tree(0)(1851); --27 bits 
            adder_tree(1)(926) <= adder_tree(0)(1852) + adder_tree(0)(1853); --27 bits 
            adder_tree(1)(927) <= adder_tree(0)(1854) + adder_tree(0)(1855); --27 bits 
            adder_tree(1)(928) <= adder_tree(0)(1856) + adder_tree(0)(1857); --27 bits 
            adder_tree(1)(929) <= adder_tree(0)(1858) + adder_tree(0)(1859); --27 bits 
            adder_tree(1)(930) <= adder_tree(0)(1860) + adder_tree(0)(1861); --27 bits 
            adder_tree(1)(931) <= adder_tree(0)(1862) + adder_tree(0)(1863); --27 bits 
            adder_tree(1)(932) <= adder_tree(0)(1864) + adder_tree(0)(1865); --27 bits 
            adder_tree(1)(933) <= adder_tree(0)(1866) + adder_tree(0)(1867); --27 bits 
            adder_tree(1)(934) <= adder_tree(0)(1868) + adder_tree(0)(1869); --27 bits 
            adder_tree(1)(935) <= adder_tree(0)(1870) + adder_tree(0)(1871); --27 bits 
            adder_tree(1)(936) <= adder_tree(0)(1872) + adder_tree(0)(1873); --27 bits 
            adder_tree(1)(937) <= adder_tree(0)(1874) + adder_tree(0)(1875); --27 bits 
            adder_tree(1)(938) <= adder_tree(0)(1876) + adder_tree(0)(1877); --27 bits 
            adder_tree(1)(939) <= adder_tree(0)(1878) + adder_tree(0)(1879); --27 bits 
            adder_tree(1)(940) <= adder_tree(0)(1880) + adder_tree(0)(1881); --27 bits 
            adder_tree(1)(941) <= adder_tree(0)(1882) + adder_tree(0)(1883); --27 bits 
            adder_tree(1)(942) <= adder_tree(0)(1884) + adder_tree(0)(1885); --27 bits 
            adder_tree(1)(943) <= adder_tree(0)(1886) + adder_tree(0)(1887); --27 bits 
            adder_tree(1)(944) <= adder_tree(0)(1888) + adder_tree(0)(1889); --27 bits 
            adder_tree(1)(945) <= adder_tree(0)(1890) + adder_tree(0)(1891); --27 bits 
            adder_tree(1)(946) <= adder_tree(0)(1892) + adder_tree(0)(1893); --27 bits 
            adder_tree(1)(947) <= adder_tree(0)(1894) + adder_tree(0)(1895); --27 bits 
            adder_tree(1)(948) <= adder_tree(0)(1896) + adder_tree(0)(1897); --27 bits 
            adder_tree(1)(949) <= adder_tree(0)(1898) + adder_tree(0)(1899); --27 bits 
            adder_tree(1)(950) <= adder_tree(0)(1900) + adder_tree(0)(1901); --27 bits 
            adder_tree(1)(951) <= adder_tree(0)(1902) + adder_tree(0)(1903); --27 bits 
            adder_tree(1)(952) <= adder_tree(0)(1904) + adder_tree(0)(1905); --27 bits 
            adder_tree(1)(953) <= adder_tree(0)(1906) + adder_tree(0)(1907); --27 bits 
            adder_tree(1)(954) <= adder_tree(0)(1908) + adder_tree(0)(1909); --27 bits 
            adder_tree(1)(955) <= adder_tree(0)(1910) + adder_tree(0)(1911); --27 bits 
            adder_tree(1)(956) <= adder_tree(0)(1912) + adder_tree(0)(1913); --27 bits 
            adder_tree(1)(957) <= adder_tree(0)(1914) + adder_tree(0)(1915); --27 bits 
            adder_tree(1)(958) <= adder_tree(0)(1916) + adder_tree(0)(1917); --27 bits 
            adder_tree(1)(959) <= adder_tree(0)(1918) + adder_tree(0)(1919); --27 bits 
            adder_tree(1)(960) <= adder_tree(0)(1920) + adder_tree(0)(1921); --27 bits 
            adder_tree(1)(961) <= adder_tree(0)(1922) + adder_tree(0)(1923); --27 bits 
            adder_tree(1)(962) <= adder_tree(0)(1924) + adder_tree(0)(1925); --27 bits 
            adder_tree(1)(963) <= adder_tree(0)(1926) + adder_tree(0)(1927); --27 bits 
            adder_tree(1)(964) <= adder_tree(0)(1928) + adder_tree(0)(1929); --27 bits 
            adder_tree(1)(965) <= adder_tree(0)(1930) + adder_tree(0)(1931); --27 bits 
            adder_tree(1)(966) <= adder_tree(0)(1932) + adder_tree(0)(1933); --27 bits 
            adder_tree(1)(967) <= adder_tree(0)(1934) + adder_tree(0)(1935); --27 bits 
            adder_tree(1)(968) <= adder_tree(0)(1936) + adder_tree(0)(1937); --27 bits 
            adder_tree(1)(969) <= adder_tree(0)(1938) + adder_tree(0)(1939); --27 bits 
            adder_tree(1)(970) <= adder_tree(0)(1940) + adder_tree(0)(1941); --27 bits 
            adder_tree(1)(971) <= adder_tree(0)(1942) + adder_tree(0)(1943); --27 bits 
            adder_tree(1)(972) <= adder_tree(0)(1944) + adder_tree(0)(1945); --27 bits 
            adder_tree(1)(973) <= adder_tree(0)(1946) + adder_tree(0)(1947); --27 bits 
            adder_tree(1)(974) <= adder_tree(0)(1948) + adder_tree(0)(1949); --27 bits 
            adder_tree(1)(975) <= adder_tree(0)(1950) + adder_tree(0)(1951); --27 bits 
            adder_tree(1)(976) <= adder_tree(0)(1952) + adder_tree(0)(1953); --27 bits 
            adder_tree(1)(977) <= adder_tree(0)(1954) + adder_tree(0)(1955); --27 bits 
            adder_tree(1)(978) <= adder_tree(0)(1956) + adder_tree(0)(1957); --27 bits 
            adder_tree(1)(979) <= adder_tree(0)(1958) + adder_tree(0)(1959); --27 bits 
            adder_tree(1)(980) <= adder_tree(0)(1960) + adder_tree(0)(1961); --27 bits 
            adder_tree(1)(981) <= adder_tree(0)(1962) + adder_tree(0)(1963); --27 bits 
            adder_tree(1)(982) <= adder_tree(0)(1964) + adder_tree(0)(1965); --27 bits 
            adder_tree(1)(983) <= adder_tree(0)(1966) + adder_tree(0)(1967); --27 bits 
            adder_tree(1)(984) <= adder_tree(0)(1968) + adder_tree(0)(1969); --27 bits 
            adder_tree(1)(985) <= adder_tree(0)(1970) + adder_tree(0)(1971); --27 bits 
            adder_tree(1)(986) <= adder_tree(0)(1972) + adder_tree(0)(1973); --27 bits 
            adder_tree(1)(987) <= adder_tree(0)(1974) + adder_tree(0)(1975); --27 bits 
            adder_tree(1)(988) <= adder_tree(0)(1976) + adder_tree(0)(1977); --27 bits 
            adder_tree(1)(989) <= adder_tree(0)(1978) + adder_tree(0)(1979); --27 bits 
            adder_tree(1)(990) <= adder_tree(0)(1980) + adder_tree(0)(1981); --27 bits 
            adder_tree(1)(991) <= adder_tree(0)(1982) + adder_tree(0)(1983); --27 bits 
            adder_tree(1)(992) <= adder_tree(0)(1984) + adder_tree(0)(1985); --27 bits 
            adder_tree(1)(993) <= adder_tree(0)(1986) + adder_tree(0)(1987); --27 bits 
            adder_tree(1)(994) <= adder_tree(0)(1988) + adder_tree(0)(1989); --27 bits 
            adder_tree(1)(995) <= adder_tree(0)(1990) + adder_tree(0)(1991); --27 bits 
            adder_tree(1)(996) <= adder_tree(0)(1992) + adder_tree(0)(1993); --27 bits 
            adder_tree(1)(997) <= adder_tree(0)(1994) + adder_tree(0)(1995); --27 bits 
            adder_tree(1)(998) <= adder_tree(0)(1996) + adder_tree(0)(1997); --27 bits 
            adder_tree(1)(999) <= adder_tree(0)(1998) + adder_tree(0)(1999); --27 bits 
            adder_tree(1)(1000) <= adder_tree(0)(2000) + adder_tree(0)(2001); --27 bits 
            adder_tree(1)(1001) <= adder_tree(0)(2002) + adder_tree(0)(2003); --27 bits 
            adder_tree(1)(1002) <= adder_tree(0)(2004) + adder_tree(0)(2005); --27 bits 
            adder_tree(1)(1003) <= adder_tree(0)(2006) + adder_tree(0)(2007); --27 bits 
            adder_tree(1)(1004) <= adder_tree(0)(2008) + adder_tree(0)(2009); --27 bits 
            adder_tree(1)(1005) <= adder_tree(0)(2010) + adder_tree(0)(2011); --27 bits 
            adder_tree(1)(1006) <= adder_tree(0)(2012) + adder_tree(0)(2013); --27 bits 
            adder_tree(1)(1007) <= adder_tree(0)(2014) + adder_tree(0)(2015); --27 bits 
            adder_tree(1)(1008) <= adder_tree(0)(2016) + adder_tree(0)(2017); --27 bits 
            adder_tree(1)(1009) <= adder_tree(0)(2018) + adder_tree(0)(2019); --27 bits 
            adder_tree(1)(1010) <= adder_tree(0)(2020) + adder_tree(0)(2021); --27 bits 
            adder_tree(1)(1011) <= adder_tree(0)(2022) + adder_tree(0)(2023); --27 bits 
            adder_tree(1)(1012) <= adder_tree(0)(2024) + adder_tree(0)(2025); --27 bits 
            adder_tree(1)(1013) <= adder_tree(0)(2026) + adder_tree(0)(2027); --27 bits 
            adder_tree(1)(1014) <= adder_tree(0)(2028) + adder_tree(0)(2029); --27 bits 
            adder_tree(1)(1015) <= adder_tree(0)(2030) + adder_tree(0)(2031); --27 bits 
            adder_tree(1)(1016) <= adder_tree(0)(2032) + adder_tree(0)(2033); --27 bits 
            adder_tree(1)(1017) <= adder_tree(0)(2034) + adder_tree(0)(2035); --27 bits 
            adder_tree(1)(1018) <= adder_tree(0)(2036) + adder_tree(0)(2037); --27 bits 
            adder_tree(1)(1019) <= adder_tree(0)(2038) + adder_tree(0)(2039); --27 bits 
            adder_tree(1)(1020) <= adder_tree(0)(2040) + adder_tree(0)(2041); --27 bits 
            adder_tree(1)(1021) <= adder_tree(0)(2042) + adder_tree(0)(2043); --27 bits 
            adder_tree(1)(1022) <= adder_tree(0)(2044) + adder_tree(0)(2045); --27 bits 
            adder_tree(1)(1023) <= adder_tree(0)(2046) + adder_tree(0)(2047); --27 bits 
            adder_tree(2)(0) <= adder_tree(1)(0) + adder_tree(1)(1); --28 bits 
            adder_tree(2)(1) <= adder_tree(1)(2) + adder_tree(1)(3); --28 bits 
            adder_tree(2)(2) <= adder_tree(1)(4) + adder_tree(1)(5); --28 bits 
            adder_tree(2)(3) <= adder_tree(1)(6) + adder_tree(1)(7); --28 bits 
            adder_tree(2)(4) <= adder_tree(1)(8) + adder_tree(1)(9); --28 bits 
            adder_tree(2)(5) <= adder_tree(1)(10) + adder_tree(1)(11); --28 bits 
            adder_tree(2)(6) <= adder_tree(1)(12) + adder_tree(1)(13); --28 bits 
            adder_tree(2)(7) <= adder_tree(1)(14) + adder_tree(1)(15); --28 bits 
            adder_tree(2)(8) <= adder_tree(1)(16) + adder_tree(1)(17); --28 bits 
            adder_tree(2)(9) <= adder_tree(1)(18) + adder_tree(1)(19); --28 bits 
            adder_tree(2)(10) <= adder_tree(1)(20) + adder_tree(1)(21); --28 bits 
            adder_tree(2)(11) <= adder_tree(1)(22) + adder_tree(1)(23); --28 bits 
            adder_tree(2)(12) <= adder_tree(1)(24) + adder_tree(1)(25); --28 bits 
            adder_tree(2)(13) <= adder_tree(1)(26) + adder_tree(1)(27); --28 bits 
            adder_tree(2)(14) <= adder_tree(1)(28) + adder_tree(1)(29); --28 bits 
            adder_tree(2)(15) <= adder_tree(1)(30) + adder_tree(1)(31); --28 bits 
            adder_tree(2)(16) <= adder_tree(1)(32) + adder_tree(1)(33); --28 bits 
            adder_tree(2)(17) <= adder_tree(1)(34) + adder_tree(1)(35); --28 bits 
            adder_tree(2)(18) <= adder_tree(1)(36) + adder_tree(1)(37); --28 bits 
            adder_tree(2)(19) <= adder_tree(1)(38) + adder_tree(1)(39); --28 bits 
            adder_tree(2)(20) <= adder_tree(1)(40) + adder_tree(1)(41); --28 bits 
            adder_tree(2)(21) <= adder_tree(1)(42) + adder_tree(1)(43); --28 bits 
            adder_tree(2)(22) <= adder_tree(1)(44) + adder_tree(1)(45); --28 bits 
            adder_tree(2)(23) <= adder_tree(1)(46) + adder_tree(1)(47); --28 bits 
            adder_tree(2)(24) <= adder_tree(1)(48) + adder_tree(1)(49); --28 bits 
            adder_tree(2)(25) <= adder_tree(1)(50) + adder_tree(1)(51); --28 bits 
            adder_tree(2)(26) <= adder_tree(1)(52) + adder_tree(1)(53); --28 bits 
            adder_tree(2)(27) <= adder_tree(1)(54) + adder_tree(1)(55); --28 bits 
            adder_tree(2)(28) <= adder_tree(1)(56) + adder_tree(1)(57); --28 bits 
            adder_tree(2)(29) <= adder_tree(1)(58) + adder_tree(1)(59); --28 bits 
            adder_tree(2)(30) <= adder_tree(1)(60) + adder_tree(1)(61); --28 bits 
            adder_tree(2)(31) <= adder_tree(1)(62) + adder_tree(1)(63); --28 bits 
            adder_tree(2)(32) <= adder_tree(1)(64) + adder_tree(1)(65); --28 bits 
            adder_tree(2)(33) <= adder_tree(1)(66) + adder_tree(1)(67); --28 bits 
            adder_tree(2)(34) <= adder_tree(1)(68) + adder_tree(1)(69); --28 bits 
            adder_tree(2)(35) <= adder_tree(1)(70) + adder_tree(1)(71); --28 bits 
            adder_tree(2)(36) <= adder_tree(1)(72) + adder_tree(1)(73); --28 bits 
            adder_tree(2)(37) <= adder_tree(1)(74) + adder_tree(1)(75); --28 bits 
            adder_tree(2)(38) <= adder_tree(1)(76) + adder_tree(1)(77); --28 bits 
            adder_tree(2)(39) <= adder_tree(1)(78) + adder_tree(1)(79); --28 bits 
            adder_tree(2)(40) <= adder_tree(1)(80) + adder_tree(1)(81); --28 bits 
            adder_tree(2)(41) <= adder_tree(1)(82) + adder_tree(1)(83); --28 bits 
            adder_tree(2)(42) <= adder_tree(1)(84) + adder_tree(1)(85); --28 bits 
            adder_tree(2)(43) <= adder_tree(1)(86) + adder_tree(1)(87); --28 bits 
            adder_tree(2)(44) <= adder_tree(1)(88) + adder_tree(1)(89); --28 bits 
            adder_tree(2)(45) <= adder_tree(1)(90) + adder_tree(1)(91); --28 bits 
            adder_tree(2)(46) <= adder_tree(1)(92) + adder_tree(1)(93); --28 bits 
            adder_tree(2)(47) <= adder_tree(1)(94) + adder_tree(1)(95); --28 bits 
            adder_tree(2)(48) <= adder_tree(1)(96) + adder_tree(1)(97); --28 bits 
            adder_tree(2)(49) <= adder_tree(1)(98) + adder_tree(1)(99); --28 bits 
            adder_tree(2)(50) <= adder_tree(1)(100) + adder_tree(1)(101); --28 bits 
            adder_tree(2)(51) <= adder_tree(1)(102) + adder_tree(1)(103); --28 bits 
            adder_tree(2)(52) <= adder_tree(1)(104) + adder_tree(1)(105); --28 bits 
            adder_tree(2)(53) <= adder_tree(1)(106) + adder_tree(1)(107); --28 bits 
            adder_tree(2)(54) <= adder_tree(1)(108) + adder_tree(1)(109); --28 bits 
            adder_tree(2)(55) <= adder_tree(1)(110) + adder_tree(1)(111); --28 bits 
            adder_tree(2)(56) <= adder_tree(1)(112) + adder_tree(1)(113); --28 bits 
            adder_tree(2)(57) <= adder_tree(1)(114) + adder_tree(1)(115); --28 bits 
            adder_tree(2)(58) <= adder_tree(1)(116) + adder_tree(1)(117); --28 bits 
            adder_tree(2)(59) <= adder_tree(1)(118) + adder_tree(1)(119); --28 bits 
            adder_tree(2)(60) <= adder_tree(1)(120) + adder_tree(1)(121); --28 bits 
            adder_tree(2)(61) <= adder_tree(1)(122) + adder_tree(1)(123); --28 bits 
            adder_tree(2)(62) <= adder_tree(1)(124) + adder_tree(1)(125); --28 bits 
            adder_tree(2)(63) <= adder_tree(1)(126) + adder_tree(1)(127); --28 bits 
            adder_tree(2)(64) <= adder_tree(1)(128) + adder_tree(1)(129); --28 bits 
            adder_tree(2)(65) <= adder_tree(1)(130) + adder_tree(1)(131); --28 bits 
            adder_tree(2)(66) <= adder_tree(1)(132) + adder_tree(1)(133); --28 bits 
            adder_tree(2)(67) <= adder_tree(1)(134) + adder_tree(1)(135); --28 bits 
            adder_tree(2)(68) <= adder_tree(1)(136) + adder_tree(1)(137); --28 bits 
            adder_tree(2)(69) <= adder_tree(1)(138) + adder_tree(1)(139); --28 bits 
            adder_tree(2)(70) <= adder_tree(1)(140) + adder_tree(1)(141); --28 bits 
            adder_tree(2)(71) <= adder_tree(1)(142) + adder_tree(1)(143); --28 bits 
            adder_tree(2)(72) <= adder_tree(1)(144) + adder_tree(1)(145); --28 bits 
            adder_tree(2)(73) <= adder_tree(1)(146) + adder_tree(1)(147); --28 bits 
            adder_tree(2)(74) <= adder_tree(1)(148) + adder_tree(1)(149); --28 bits 
            adder_tree(2)(75) <= adder_tree(1)(150) + adder_tree(1)(151); --28 bits 
            adder_tree(2)(76) <= adder_tree(1)(152) + adder_tree(1)(153); --28 bits 
            adder_tree(2)(77) <= adder_tree(1)(154) + adder_tree(1)(155); --28 bits 
            adder_tree(2)(78) <= adder_tree(1)(156) + adder_tree(1)(157); --28 bits 
            adder_tree(2)(79) <= adder_tree(1)(158) + adder_tree(1)(159); --28 bits 
            adder_tree(2)(80) <= adder_tree(1)(160) + adder_tree(1)(161); --28 bits 
            adder_tree(2)(81) <= adder_tree(1)(162) + adder_tree(1)(163); --28 bits 
            adder_tree(2)(82) <= adder_tree(1)(164) + adder_tree(1)(165); --28 bits 
            adder_tree(2)(83) <= adder_tree(1)(166) + adder_tree(1)(167); --28 bits 
            adder_tree(2)(84) <= adder_tree(1)(168) + adder_tree(1)(169); --28 bits 
            adder_tree(2)(85) <= adder_tree(1)(170) + adder_tree(1)(171); --28 bits 
            adder_tree(2)(86) <= adder_tree(1)(172) + adder_tree(1)(173); --28 bits 
            adder_tree(2)(87) <= adder_tree(1)(174) + adder_tree(1)(175); --28 bits 
            adder_tree(2)(88) <= adder_tree(1)(176) + adder_tree(1)(177); --28 bits 
            adder_tree(2)(89) <= adder_tree(1)(178) + adder_tree(1)(179); --28 bits 
            adder_tree(2)(90) <= adder_tree(1)(180) + adder_tree(1)(181); --28 bits 
            adder_tree(2)(91) <= adder_tree(1)(182) + adder_tree(1)(183); --28 bits 
            adder_tree(2)(92) <= adder_tree(1)(184) + adder_tree(1)(185); --28 bits 
            adder_tree(2)(93) <= adder_tree(1)(186) + adder_tree(1)(187); --28 bits 
            adder_tree(2)(94) <= adder_tree(1)(188) + adder_tree(1)(189); --28 bits 
            adder_tree(2)(95) <= adder_tree(1)(190) + adder_tree(1)(191); --28 bits 
            adder_tree(2)(96) <= adder_tree(1)(192) + adder_tree(1)(193); --28 bits 
            adder_tree(2)(97) <= adder_tree(1)(194) + adder_tree(1)(195); --28 bits 
            adder_tree(2)(98) <= adder_tree(1)(196) + adder_tree(1)(197); --28 bits 
            adder_tree(2)(99) <= adder_tree(1)(198) + adder_tree(1)(199); --28 bits 
            adder_tree(2)(100) <= adder_tree(1)(200) + adder_tree(1)(201); --28 bits 
            adder_tree(2)(101) <= adder_tree(1)(202) + adder_tree(1)(203); --28 bits 
            adder_tree(2)(102) <= adder_tree(1)(204) + adder_tree(1)(205); --28 bits 
            adder_tree(2)(103) <= adder_tree(1)(206) + adder_tree(1)(207); --28 bits 
            adder_tree(2)(104) <= adder_tree(1)(208) + adder_tree(1)(209); --28 bits 
            adder_tree(2)(105) <= adder_tree(1)(210) + adder_tree(1)(211); --28 bits 
            adder_tree(2)(106) <= adder_tree(1)(212) + adder_tree(1)(213); --28 bits 
            adder_tree(2)(107) <= adder_tree(1)(214) + adder_tree(1)(215); --28 bits 
            adder_tree(2)(108) <= adder_tree(1)(216) + adder_tree(1)(217); --28 bits 
            adder_tree(2)(109) <= adder_tree(1)(218) + adder_tree(1)(219); --28 bits 
            adder_tree(2)(110) <= adder_tree(1)(220) + adder_tree(1)(221); --28 bits 
            adder_tree(2)(111) <= adder_tree(1)(222) + adder_tree(1)(223); --28 bits 
            adder_tree(2)(112) <= adder_tree(1)(224) + adder_tree(1)(225); --28 bits 
            adder_tree(2)(113) <= adder_tree(1)(226) + adder_tree(1)(227); --28 bits 
            adder_tree(2)(114) <= adder_tree(1)(228) + adder_tree(1)(229); --28 bits 
            adder_tree(2)(115) <= adder_tree(1)(230) + adder_tree(1)(231); --28 bits 
            adder_tree(2)(116) <= adder_tree(1)(232) + adder_tree(1)(233); --28 bits 
            adder_tree(2)(117) <= adder_tree(1)(234) + adder_tree(1)(235); --28 bits 
            adder_tree(2)(118) <= adder_tree(1)(236) + adder_tree(1)(237); --28 bits 
            adder_tree(2)(119) <= adder_tree(1)(238) + adder_tree(1)(239); --28 bits 
            adder_tree(2)(120) <= adder_tree(1)(240) + adder_tree(1)(241); --28 bits 
            adder_tree(2)(121) <= adder_tree(1)(242) + adder_tree(1)(243); --28 bits 
            adder_tree(2)(122) <= adder_tree(1)(244) + adder_tree(1)(245); --28 bits 
            adder_tree(2)(123) <= adder_tree(1)(246) + adder_tree(1)(247); --28 bits 
            adder_tree(2)(124) <= adder_tree(1)(248) + adder_tree(1)(249); --28 bits 
            adder_tree(2)(125) <= adder_tree(1)(250) + adder_tree(1)(251); --28 bits 
            adder_tree(2)(126) <= adder_tree(1)(252) + adder_tree(1)(253); --28 bits 
            adder_tree(2)(127) <= adder_tree(1)(254) + adder_tree(1)(255); --28 bits 
            adder_tree(2)(128) <= adder_tree(1)(256) + adder_tree(1)(257); --28 bits 
            adder_tree(2)(129) <= adder_tree(1)(258) + adder_tree(1)(259); --28 bits 
            adder_tree(2)(130) <= adder_tree(1)(260) + adder_tree(1)(261); --28 bits 
            adder_tree(2)(131) <= adder_tree(1)(262) + adder_tree(1)(263); --28 bits 
            adder_tree(2)(132) <= adder_tree(1)(264) + adder_tree(1)(265); --28 bits 
            adder_tree(2)(133) <= adder_tree(1)(266) + adder_tree(1)(267); --28 bits 
            adder_tree(2)(134) <= adder_tree(1)(268) + adder_tree(1)(269); --28 bits 
            adder_tree(2)(135) <= adder_tree(1)(270) + adder_tree(1)(271); --28 bits 
            adder_tree(2)(136) <= adder_tree(1)(272) + adder_tree(1)(273); --28 bits 
            adder_tree(2)(137) <= adder_tree(1)(274) + adder_tree(1)(275); --28 bits 
            adder_tree(2)(138) <= adder_tree(1)(276) + adder_tree(1)(277); --28 bits 
            adder_tree(2)(139) <= adder_tree(1)(278) + adder_tree(1)(279); --28 bits 
            adder_tree(2)(140) <= adder_tree(1)(280) + adder_tree(1)(281); --28 bits 
            adder_tree(2)(141) <= adder_tree(1)(282) + adder_tree(1)(283); --28 bits 
            adder_tree(2)(142) <= adder_tree(1)(284) + adder_tree(1)(285); --28 bits 
            adder_tree(2)(143) <= adder_tree(1)(286) + adder_tree(1)(287); --28 bits 
            adder_tree(2)(144) <= adder_tree(1)(288) + adder_tree(1)(289); --28 bits 
            adder_tree(2)(145) <= adder_tree(1)(290) + adder_tree(1)(291); --28 bits 
            adder_tree(2)(146) <= adder_tree(1)(292) + adder_tree(1)(293); --28 bits 
            adder_tree(2)(147) <= adder_tree(1)(294) + adder_tree(1)(295); --28 bits 
            adder_tree(2)(148) <= adder_tree(1)(296) + adder_tree(1)(297); --28 bits 
            adder_tree(2)(149) <= adder_tree(1)(298) + adder_tree(1)(299); --28 bits 
            adder_tree(2)(150) <= adder_tree(1)(300) + adder_tree(1)(301); --28 bits 
            adder_tree(2)(151) <= adder_tree(1)(302) + adder_tree(1)(303); --28 bits 
            adder_tree(2)(152) <= adder_tree(1)(304) + adder_tree(1)(305); --28 bits 
            adder_tree(2)(153) <= adder_tree(1)(306) + adder_tree(1)(307); --28 bits 
            adder_tree(2)(154) <= adder_tree(1)(308) + adder_tree(1)(309); --28 bits 
            adder_tree(2)(155) <= adder_tree(1)(310) + adder_tree(1)(311); --28 bits 
            adder_tree(2)(156) <= adder_tree(1)(312) + adder_tree(1)(313); --28 bits 
            adder_tree(2)(157) <= adder_tree(1)(314) + adder_tree(1)(315); --28 bits 
            adder_tree(2)(158) <= adder_tree(1)(316) + adder_tree(1)(317); --28 bits 
            adder_tree(2)(159) <= adder_tree(1)(318) + adder_tree(1)(319); --28 bits 
            adder_tree(2)(160) <= adder_tree(1)(320) + adder_tree(1)(321); --28 bits 
            adder_tree(2)(161) <= adder_tree(1)(322) + adder_tree(1)(323); --28 bits 
            adder_tree(2)(162) <= adder_tree(1)(324) + adder_tree(1)(325); --28 bits 
            adder_tree(2)(163) <= adder_tree(1)(326) + adder_tree(1)(327); --28 bits 
            adder_tree(2)(164) <= adder_tree(1)(328) + adder_tree(1)(329); --28 bits 
            adder_tree(2)(165) <= adder_tree(1)(330) + adder_tree(1)(331); --28 bits 
            adder_tree(2)(166) <= adder_tree(1)(332) + adder_tree(1)(333); --28 bits 
            adder_tree(2)(167) <= adder_tree(1)(334) + adder_tree(1)(335); --28 bits 
            adder_tree(2)(168) <= adder_tree(1)(336) + adder_tree(1)(337); --28 bits 
            adder_tree(2)(169) <= adder_tree(1)(338) + adder_tree(1)(339); --28 bits 
            adder_tree(2)(170) <= adder_tree(1)(340) + adder_tree(1)(341); --28 bits 
            adder_tree(2)(171) <= adder_tree(1)(342) + adder_tree(1)(343); --28 bits 
            adder_tree(2)(172) <= adder_tree(1)(344) + adder_tree(1)(345); --28 bits 
            adder_tree(2)(173) <= adder_tree(1)(346) + adder_tree(1)(347); --28 bits 
            adder_tree(2)(174) <= adder_tree(1)(348) + adder_tree(1)(349); --28 bits 
            adder_tree(2)(175) <= adder_tree(1)(350) + adder_tree(1)(351); --28 bits 
            adder_tree(2)(176) <= adder_tree(1)(352) + adder_tree(1)(353); --28 bits 
            adder_tree(2)(177) <= adder_tree(1)(354) + adder_tree(1)(355); --28 bits 
            adder_tree(2)(178) <= adder_tree(1)(356) + adder_tree(1)(357); --28 bits 
            adder_tree(2)(179) <= adder_tree(1)(358) + adder_tree(1)(359); --28 bits 
            adder_tree(2)(180) <= adder_tree(1)(360) + adder_tree(1)(361); --28 bits 
            adder_tree(2)(181) <= adder_tree(1)(362) + adder_tree(1)(363); --28 bits 
            adder_tree(2)(182) <= adder_tree(1)(364) + adder_tree(1)(365); --28 bits 
            adder_tree(2)(183) <= adder_tree(1)(366) + adder_tree(1)(367); --28 bits 
            adder_tree(2)(184) <= adder_tree(1)(368) + adder_tree(1)(369); --28 bits 
            adder_tree(2)(185) <= adder_tree(1)(370) + adder_tree(1)(371); --28 bits 
            adder_tree(2)(186) <= adder_tree(1)(372) + adder_tree(1)(373); --28 bits 
            adder_tree(2)(187) <= adder_tree(1)(374) + adder_tree(1)(375); --28 bits 
            adder_tree(2)(188) <= adder_tree(1)(376) + adder_tree(1)(377); --28 bits 
            adder_tree(2)(189) <= adder_tree(1)(378) + adder_tree(1)(379); --28 bits 
            adder_tree(2)(190) <= adder_tree(1)(380) + adder_tree(1)(381); --28 bits 
            adder_tree(2)(191) <= adder_tree(1)(382) + adder_tree(1)(383); --28 bits 
            adder_tree(2)(192) <= adder_tree(1)(384) + adder_tree(1)(385); --28 bits 
            adder_tree(2)(193) <= adder_tree(1)(386) + adder_tree(1)(387); --28 bits 
            adder_tree(2)(194) <= adder_tree(1)(388) + adder_tree(1)(389); --28 bits 
            adder_tree(2)(195) <= adder_tree(1)(390) + adder_tree(1)(391); --28 bits 
            adder_tree(2)(196) <= adder_tree(1)(392) + adder_tree(1)(393); --28 bits 
            adder_tree(2)(197) <= adder_tree(1)(394) + adder_tree(1)(395); --28 bits 
            adder_tree(2)(198) <= adder_tree(1)(396) + adder_tree(1)(397); --28 bits 
            adder_tree(2)(199) <= adder_tree(1)(398) + adder_tree(1)(399); --28 bits 
            adder_tree(2)(200) <= adder_tree(1)(400) + adder_tree(1)(401); --28 bits 
            adder_tree(2)(201) <= adder_tree(1)(402) + adder_tree(1)(403); --28 bits 
            adder_tree(2)(202) <= adder_tree(1)(404) + adder_tree(1)(405); --28 bits 
            adder_tree(2)(203) <= adder_tree(1)(406) + adder_tree(1)(407); --28 bits 
            adder_tree(2)(204) <= adder_tree(1)(408) + adder_tree(1)(409); --28 bits 
            adder_tree(2)(205) <= adder_tree(1)(410) + adder_tree(1)(411); --28 bits 
            adder_tree(2)(206) <= adder_tree(1)(412) + adder_tree(1)(413); --28 bits 
            adder_tree(2)(207) <= adder_tree(1)(414) + adder_tree(1)(415); --28 bits 
            adder_tree(2)(208) <= adder_tree(1)(416) + adder_tree(1)(417); --28 bits 
            adder_tree(2)(209) <= adder_tree(1)(418) + adder_tree(1)(419); --28 bits 
            adder_tree(2)(210) <= adder_tree(1)(420) + adder_tree(1)(421); --28 bits 
            adder_tree(2)(211) <= adder_tree(1)(422) + adder_tree(1)(423); --28 bits 
            adder_tree(2)(212) <= adder_tree(1)(424) + adder_tree(1)(425); --28 bits 
            adder_tree(2)(213) <= adder_tree(1)(426) + adder_tree(1)(427); --28 bits 
            adder_tree(2)(214) <= adder_tree(1)(428) + adder_tree(1)(429); --28 bits 
            adder_tree(2)(215) <= adder_tree(1)(430) + adder_tree(1)(431); --28 bits 
            adder_tree(2)(216) <= adder_tree(1)(432) + adder_tree(1)(433); --28 bits 
            adder_tree(2)(217) <= adder_tree(1)(434) + adder_tree(1)(435); --28 bits 
            adder_tree(2)(218) <= adder_tree(1)(436) + adder_tree(1)(437); --28 bits 
            adder_tree(2)(219) <= adder_tree(1)(438) + adder_tree(1)(439); --28 bits 
            adder_tree(2)(220) <= adder_tree(1)(440) + adder_tree(1)(441); --28 bits 
            adder_tree(2)(221) <= adder_tree(1)(442) + adder_tree(1)(443); --28 bits 
            adder_tree(2)(222) <= adder_tree(1)(444) + adder_tree(1)(445); --28 bits 
            adder_tree(2)(223) <= adder_tree(1)(446) + adder_tree(1)(447); --28 bits 
            adder_tree(2)(224) <= adder_tree(1)(448) + adder_tree(1)(449); --28 bits 
            adder_tree(2)(225) <= adder_tree(1)(450) + adder_tree(1)(451); --28 bits 
            adder_tree(2)(226) <= adder_tree(1)(452) + adder_tree(1)(453); --28 bits 
            adder_tree(2)(227) <= adder_tree(1)(454) + adder_tree(1)(455); --28 bits 
            adder_tree(2)(228) <= adder_tree(1)(456) + adder_tree(1)(457); --28 bits 
            adder_tree(2)(229) <= adder_tree(1)(458) + adder_tree(1)(459); --28 bits 
            adder_tree(2)(230) <= adder_tree(1)(460) + adder_tree(1)(461); --28 bits 
            adder_tree(2)(231) <= adder_tree(1)(462) + adder_tree(1)(463); --28 bits 
            adder_tree(2)(232) <= adder_tree(1)(464) + adder_tree(1)(465); --28 bits 
            adder_tree(2)(233) <= adder_tree(1)(466) + adder_tree(1)(467); --28 bits 
            adder_tree(2)(234) <= adder_tree(1)(468) + adder_tree(1)(469); --28 bits 
            adder_tree(2)(235) <= adder_tree(1)(470) + adder_tree(1)(471); --28 bits 
            adder_tree(2)(236) <= adder_tree(1)(472) + adder_tree(1)(473); --28 bits 
            adder_tree(2)(237) <= adder_tree(1)(474) + adder_tree(1)(475); --28 bits 
            adder_tree(2)(238) <= adder_tree(1)(476) + adder_tree(1)(477); --28 bits 
            adder_tree(2)(239) <= adder_tree(1)(478) + adder_tree(1)(479); --28 bits 
            adder_tree(2)(240) <= adder_tree(1)(480) + adder_tree(1)(481); --28 bits 
            adder_tree(2)(241) <= adder_tree(1)(482) + adder_tree(1)(483); --28 bits 
            adder_tree(2)(242) <= adder_tree(1)(484) + adder_tree(1)(485); --28 bits 
            adder_tree(2)(243) <= adder_tree(1)(486) + adder_tree(1)(487); --28 bits 
            adder_tree(2)(244) <= adder_tree(1)(488) + adder_tree(1)(489); --28 bits 
            adder_tree(2)(245) <= adder_tree(1)(490) + adder_tree(1)(491); --28 bits 
            adder_tree(2)(246) <= adder_tree(1)(492) + adder_tree(1)(493); --28 bits 
            adder_tree(2)(247) <= adder_tree(1)(494) + adder_tree(1)(495); --28 bits 
            adder_tree(2)(248) <= adder_tree(1)(496) + adder_tree(1)(497); --28 bits 
            adder_tree(2)(249) <= adder_tree(1)(498) + adder_tree(1)(499); --28 bits 
            adder_tree(2)(250) <= adder_tree(1)(500) + adder_tree(1)(501); --28 bits 
            adder_tree(2)(251) <= adder_tree(1)(502) + adder_tree(1)(503); --28 bits 
            adder_tree(2)(252) <= adder_tree(1)(504) + adder_tree(1)(505); --28 bits 
            adder_tree(2)(253) <= adder_tree(1)(506) + adder_tree(1)(507); --28 bits 
            adder_tree(2)(254) <= adder_tree(1)(508) + adder_tree(1)(509); --28 bits 
            adder_tree(2)(255) <= adder_tree(1)(510) + adder_tree(1)(511); --28 bits 
            adder_tree(2)(256) <= adder_tree(1)(512) + adder_tree(1)(513); --28 bits 
            adder_tree(2)(257) <= adder_tree(1)(514) + adder_tree(1)(515); --28 bits 
            adder_tree(2)(258) <= adder_tree(1)(516) + adder_tree(1)(517); --28 bits 
            adder_tree(2)(259) <= adder_tree(1)(518) + adder_tree(1)(519); --28 bits 
            adder_tree(2)(260) <= adder_tree(1)(520) + adder_tree(1)(521); --28 bits 
            adder_tree(2)(261) <= adder_tree(1)(522) + adder_tree(1)(523); --28 bits 
            adder_tree(2)(262) <= adder_tree(1)(524) + adder_tree(1)(525); --28 bits 
            adder_tree(2)(263) <= adder_tree(1)(526) + adder_tree(1)(527); --28 bits 
            adder_tree(2)(264) <= adder_tree(1)(528) + adder_tree(1)(529); --28 bits 
            adder_tree(2)(265) <= adder_tree(1)(530) + adder_tree(1)(531); --28 bits 
            adder_tree(2)(266) <= adder_tree(1)(532) + adder_tree(1)(533); --28 bits 
            adder_tree(2)(267) <= adder_tree(1)(534) + adder_tree(1)(535); --28 bits 
            adder_tree(2)(268) <= adder_tree(1)(536) + adder_tree(1)(537); --28 bits 
            adder_tree(2)(269) <= adder_tree(1)(538) + adder_tree(1)(539); --28 bits 
            adder_tree(2)(270) <= adder_tree(1)(540) + adder_tree(1)(541); --28 bits 
            adder_tree(2)(271) <= adder_tree(1)(542) + adder_tree(1)(543); --28 bits 
            adder_tree(2)(272) <= adder_tree(1)(544) + adder_tree(1)(545); --28 bits 
            adder_tree(2)(273) <= adder_tree(1)(546) + adder_tree(1)(547); --28 bits 
            adder_tree(2)(274) <= adder_tree(1)(548) + adder_tree(1)(549); --28 bits 
            adder_tree(2)(275) <= adder_tree(1)(550) + adder_tree(1)(551); --28 bits 
            adder_tree(2)(276) <= adder_tree(1)(552) + adder_tree(1)(553); --28 bits 
            adder_tree(2)(277) <= adder_tree(1)(554) + adder_tree(1)(555); --28 bits 
            adder_tree(2)(278) <= adder_tree(1)(556) + adder_tree(1)(557); --28 bits 
            adder_tree(2)(279) <= adder_tree(1)(558) + adder_tree(1)(559); --28 bits 
            adder_tree(2)(280) <= adder_tree(1)(560) + adder_tree(1)(561); --28 bits 
            adder_tree(2)(281) <= adder_tree(1)(562) + adder_tree(1)(563); --28 bits 
            adder_tree(2)(282) <= adder_tree(1)(564) + adder_tree(1)(565); --28 bits 
            adder_tree(2)(283) <= adder_tree(1)(566) + adder_tree(1)(567); --28 bits 
            adder_tree(2)(284) <= adder_tree(1)(568) + adder_tree(1)(569); --28 bits 
            adder_tree(2)(285) <= adder_tree(1)(570) + adder_tree(1)(571); --28 bits 
            adder_tree(2)(286) <= adder_tree(1)(572) + adder_tree(1)(573); --28 bits 
            adder_tree(2)(287) <= adder_tree(1)(574) + adder_tree(1)(575); --28 bits 
            adder_tree(2)(288) <= adder_tree(1)(576) + adder_tree(1)(577); --28 bits 
            adder_tree(2)(289) <= adder_tree(1)(578) + adder_tree(1)(579); --28 bits 
            adder_tree(2)(290) <= adder_tree(1)(580) + adder_tree(1)(581); --28 bits 
            adder_tree(2)(291) <= adder_tree(1)(582) + adder_tree(1)(583); --28 bits 
            adder_tree(2)(292) <= adder_tree(1)(584) + adder_tree(1)(585); --28 bits 
            adder_tree(2)(293) <= adder_tree(1)(586) + adder_tree(1)(587); --28 bits 
            adder_tree(2)(294) <= adder_tree(1)(588) + adder_tree(1)(589); --28 bits 
            adder_tree(2)(295) <= adder_tree(1)(590) + adder_tree(1)(591); --28 bits 
            adder_tree(2)(296) <= adder_tree(1)(592) + adder_tree(1)(593); --28 bits 
            adder_tree(2)(297) <= adder_tree(1)(594) + adder_tree(1)(595); --28 bits 
            adder_tree(2)(298) <= adder_tree(1)(596) + adder_tree(1)(597); --28 bits 
            adder_tree(2)(299) <= adder_tree(1)(598) + adder_tree(1)(599); --28 bits 
            adder_tree(2)(300) <= adder_tree(1)(600) + adder_tree(1)(601); --28 bits 
            adder_tree(2)(301) <= adder_tree(1)(602) + adder_tree(1)(603); --28 bits 
            adder_tree(2)(302) <= adder_tree(1)(604) + adder_tree(1)(605); --28 bits 
            adder_tree(2)(303) <= adder_tree(1)(606) + adder_tree(1)(607); --28 bits 
            adder_tree(2)(304) <= adder_tree(1)(608) + adder_tree(1)(609); --28 bits 
            adder_tree(2)(305) <= adder_tree(1)(610) + adder_tree(1)(611); --28 bits 
            adder_tree(2)(306) <= adder_tree(1)(612) + adder_tree(1)(613); --28 bits 
            adder_tree(2)(307) <= adder_tree(1)(614) + adder_tree(1)(615); --28 bits 
            adder_tree(2)(308) <= adder_tree(1)(616) + adder_tree(1)(617); --28 bits 
            adder_tree(2)(309) <= adder_tree(1)(618) + adder_tree(1)(619); --28 bits 
            adder_tree(2)(310) <= adder_tree(1)(620) + adder_tree(1)(621); --28 bits 
            adder_tree(2)(311) <= adder_tree(1)(622) + adder_tree(1)(623); --28 bits 
            adder_tree(2)(312) <= adder_tree(1)(624) + adder_tree(1)(625); --28 bits 
            adder_tree(2)(313) <= adder_tree(1)(626) + adder_tree(1)(627); --28 bits 
            adder_tree(2)(314) <= adder_tree(1)(628) + adder_tree(1)(629); --28 bits 
            adder_tree(2)(315) <= adder_tree(1)(630) + adder_tree(1)(631); --28 bits 
            adder_tree(2)(316) <= adder_tree(1)(632) + adder_tree(1)(633); --28 bits 
            adder_tree(2)(317) <= adder_tree(1)(634) + adder_tree(1)(635); --28 bits 
            adder_tree(2)(318) <= adder_tree(1)(636) + adder_tree(1)(637); --28 bits 
            adder_tree(2)(319) <= adder_tree(1)(638) + adder_tree(1)(639); --28 bits 
            adder_tree(2)(320) <= adder_tree(1)(640) + adder_tree(1)(641); --28 bits 
            adder_tree(2)(321) <= adder_tree(1)(642) + adder_tree(1)(643); --28 bits 
            adder_tree(2)(322) <= adder_tree(1)(644) + adder_tree(1)(645); --28 bits 
            adder_tree(2)(323) <= adder_tree(1)(646) + adder_tree(1)(647); --28 bits 
            adder_tree(2)(324) <= adder_tree(1)(648) + adder_tree(1)(649); --28 bits 
            adder_tree(2)(325) <= adder_tree(1)(650) + adder_tree(1)(651); --28 bits 
            adder_tree(2)(326) <= adder_tree(1)(652) + adder_tree(1)(653); --28 bits 
            adder_tree(2)(327) <= adder_tree(1)(654) + adder_tree(1)(655); --28 bits 
            adder_tree(2)(328) <= adder_tree(1)(656) + adder_tree(1)(657); --28 bits 
            adder_tree(2)(329) <= adder_tree(1)(658) + adder_tree(1)(659); --28 bits 
            adder_tree(2)(330) <= adder_tree(1)(660) + adder_tree(1)(661); --28 bits 
            adder_tree(2)(331) <= adder_tree(1)(662) + adder_tree(1)(663); --28 bits 
            adder_tree(2)(332) <= adder_tree(1)(664) + adder_tree(1)(665); --28 bits 
            adder_tree(2)(333) <= adder_tree(1)(666) + adder_tree(1)(667); --28 bits 
            adder_tree(2)(334) <= adder_tree(1)(668) + adder_tree(1)(669); --28 bits 
            adder_tree(2)(335) <= adder_tree(1)(670) + adder_tree(1)(671); --28 bits 
            adder_tree(2)(336) <= adder_tree(1)(672) + adder_tree(1)(673); --28 bits 
            adder_tree(2)(337) <= adder_tree(1)(674) + adder_tree(1)(675); --28 bits 
            adder_tree(2)(338) <= adder_tree(1)(676) + adder_tree(1)(677); --28 bits 
            adder_tree(2)(339) <= adder_tree(1)(678) + adder_tree(1)(679); --28 bits 
            adder_tree(2)(340) <= adder_tree(1)(680) + adder_tree(1)(681); --28 bits 
            adder_tree(2)(341) <= adder_tree(1)(682) + adder_tree(1)(683); --28 bits 
            adder_tree(2)(342) <= adder_tree(1)(684) + adder_tree(1)(685); --28 bits 
            adder_tree(2)(343) <= adder_tree(1)(686) + adder_tree(1)(687); --28 bits 
            adder_tree(2)(344) <= adder_tree(1)(688) + adder_tree(1)(689); --28 bits 
            adder_tree(2)(345) <= adder_tree(1)(690) + adder_tree(1)(691); --28 bits 
            adder_tree(2)(346) <= adder_tree(1)(692) + adder_tree(1)(693); --28 bits 
            adder_tree(2)(347) <= adder_tree(1)(694) + adder_tree(1)(695); --28 bits 
            adder_tree(2)(348) <= adder_tree(1)(696) + adder_tree(1)(697); --28 bits 
            adder_tree(2)(349) <= adder_tree(1)(698) + adder_tree(1)(699); --28 bits 
            adder_tree(2)(350) <= adder_tree(1)(700) + adder_tree(1)(701); --28 bits 
            adder_tree(2)(351) <= adder_tree(1)(702) + adder_tree(1)(703); --28 bits 
            adder_tree(2)(352) <= adder_tree(1)(704) + adder_tree(1)(705); --28 bits 
            adder_tree(2)(353) <= adder_tree(1)(706) + adder_tree(1)(707); --28 bits 
            adder_tree(2)(354) <= adder_tree(1)(708) + adder_tree(1)(709); --28 bits 
            adder_tree(2)(355) <= adder_tree(1)(710) + adder_tree(1)(711); --28 bits 
            adder_tree(2)(356) <= adder_tree(1)(712) + adder_tree(1)(713); --28 bits 
            adder_tree(2)(357) <= adder_tree(1)(714) + adder_tree(1)(715); --28 bits 
            adder_tree(2)(358) <= adder_tree(1)(716) + adder_tree(1)(717); --28 bits 
            adder_tree(2)(359) <= adder_tree(1)(718) + adder_tree(1)(719); --28 bits 
            adder_tree(2)(360) <= adder_tree(1)(720) + adder_tree(1)(721); --28 bits 
            adder_tree(2)(361) <= adder_tree(1)(722) + adder_tree(1)(723); --28 bits 
            adder_tree(2)(362) <= adder_tree(1)(724) + adder_tree(1)(725); --28 bits 
            adder_tree(2)(363) <= adder_tree(1)(726) + adder_tree(1)(727); --28 bits 
            adder_tree(2)(364) <= adder_tree(1)(728) + adder_tree(1)(729); --28 bits 
            adder_tree(2)(365) <= adder_tree(1)(730) + adder_tree(1)(731); --28 bits 
            adder_tree(2)(366) <= adder_tree(1)(732) + adder_tree(1)(733); --28 bits 
            adder_tree(2)(367) <= adder_tree(1)(734) + adder_tree(1)(735); --28 bits 
            adder_tree(2)(368) <= adder_tree(1)(736) + adder_tree(1)(737); --28 bits 
            adder_tree(2)(369) <= adder_tree(1)(738) + adder_tree(1)(739); --28 bits 
            adder_tree(2)(370) <= adder_tree(1)(740) + adder_tree(1)(741); --28 bits 
            adder_tree(2)(371) <= adder_tree(1)(742) + adder_tree(1)(743); --28 bits 
            adder_tree(2)(372) <= adder_tree(1)(744) + adder_tree(1)(745); --28 bits 
            adder_tree(2)(373) <= adder_tree(1)(746) + adder_tree(1)(747); --28 bits 
            adder_tree(2)(374) <= adder_tree(1)(748) + adder_tree(1)(749); --28 bits 
            adder_tree(2)(375) <= adder_tree(1)(750) + adder_tree(1)(751); --28 bits 
            adder_tree(2)(376) <= adder_tree(1)(752) + adder_tree(1)(753); --28 bits 
            adder_tree(2)(377) <= adder_tree(1)(754) + adder_tree(1)(755); --28 bits 
            adder_tree(2)(378) <= adder_tree(1)(756) + adder_tree(1)(757); --28 bits 
            adder_tree(2)(379) <= adder_tree(1)(758) + adder_tree(1)(759); --28 bits 
            adder_tree(2)(380) <= adder_tree(1)(760) + adder_tree(1)(761); --28 bits 
            adder_tree(2)(381) <= adder_tree(1)(762) + adder_tree(1)(763); --28 bits 
            adder_tree(2)(382) <= adder_tree(1)(764) + adder_tree(1)(765); --28 bits 
            adder_tree(2)(383) <= adder_tree(1)(766) + adder_tree(1)(767); --28 bits 
            adder_tree(2)(384) <= adder_tree(1)(768) + adder_tree(1)(769); --28 bits 
            adder_tree(2)(385) <= adder_tree(1)(770) + adder_tree(1)(771); --28 bits 
            adder_tree(2)(386) <= adder_tree(1)(772) + adder_tree(1)(773); --28 bits 
            adder_tree(2)(387) <= adder_tree(1)(774) + adder_tree(1)(775); --28 bits 
            adder_tree(2)(388) <= adder_tree(1)(776) + adder_tree(1)(777); --28 bits 
            adder_tree(2)(389) <= adder_tree(1)(778) + adder_tree(1)(779); --28 bits 
            adder_tree(2)(390) <= adder_tree(1)(780) + adder_tree(1)(781); --28 bits 
            adder_tree(2)(391) <= adder_tree(1)(782) + adder_tree(1)(783); --28 bits 
            adder_tree(2)(392) <= adder_tree(1)(784) + adder_tree(1)(785); --28 bits 
            adder_tree(2)(393) <= adder_tree(1)(786) + adder_tree(1)(787); --28 bits 
            adder_tree(2)(394) <= adder_tree(1)(788) + adder_tree(1)(789); --28 bits 
            adder_tree(2)(395) <= adder_tree(1)(790) + adder_tree(1)(791); --28 bits 
            adder_tree(2)(396) <= adder_tree(1)(792) + adder_tree(1)(793); --28 bits 
            adder_tree(2)(397) <= adder_tree(1)(794) + adder_tree(1)(795); --28 bits 
            adder_tree(2)(398) <= adder_tree(1)(796) + adder_tree(1)(797); --28 bits 
            adder_tree(2)(399) <= adder_tree(1)(798) + adder_tree(1)(799); --28 bits 
            adder_tree(2)(400) <= adder_tree(1)(800) + adder_tree(1)(801); --28 bits 
            adder_tree(2)(401) <= adder_tree(1)(802) + adder_tree(1)(803); --28 bits 
            adder_tree(2)(402) <= adder_tree(1)(804) + adder_tree(1)(805); --28 bits 
            adder_tree(2)(403) <= adder_tree(1)(806) + adder_tree(1)(807); --28 bits 
            adder_tree(2)(404) <= adder_tree(1)(808) + adder_tree(1)(809); --28 bits 
            adder_tree(2)(405) <= adder_tree(1)(810) + adder_tree(1)(811); --28 bits 
            adder_tree(2)(406) <= adder_tree(1)(812) + adder_tree(1)(813); --28 bits 
            adder_tree(2)(407) <= adder_tree(1)(814) + adder_tree(1)(815); --28 bits 
            adder_tree(2)(408) <= adder_tree(1)(816) + adder_tree(1)(817); --28 bits 
            adder_tree(2)(409) <= adder_tree(1)(818) + adder_tree(1)(819); --28 bits 
            adder_tree(2)(410) <= adder_tree(1)(820) + adder_tree(1)(821); --28 bits 
            adder_tree(2)(411) <= adder_tree(1)(822) + adder_tree(1)(823); --28 bits 
            adder_tree(2)(412) <= adder_tree(1)(824) + adder_tree(1)(825); --28 bits 
            adder_tree(2)(413) <= adder_tree(1)(826) + adder_tree(1)(827); --28 bits 
            adder_tree(2)(414) <= adder_tree(1)(828) + adder_tree(1)(829); --28 bits 
            adder_tree(2)(415) <= adder_tree(1)(830) + adder_tree(1)(831); --28 bits 
            adder_tree(2)(416) <= adder_tree(1)(832) + adder_tree(1)(833); --28 bits 
            adder_tree(2)(417) <= adder_tree(1)(834) + adder_tree(1)(835); --28 bits 
            adder_tree(2)(418) <= adder_tree(1)(836) + adder_tree(1)(837); --28 bits 
            adder_tree(2)(419) <= adder_tree(1)(838) + adder_tree(1)(839); --28 bits 
            adder_tree(2)(420) <= adder_tree(1)(840) + adder_tree(1)(841); --28 bits 
            adder_tree(2)(421) <= adder_tree(1)(842) + adder_tree(1)(843); --28 bits 
            adder_tree(2)(422) <= adder_tree(1)(844) + adder_tree(1)(845); --28 bits 
            adder_tree(2)(423) <= adder_tree(1)(846) + adder_tree(1)(847); --28 bits 
            adder_tree(2)(424) <= adder_tree(1)(848) + adder_tree(1)(849); --28 bits 
            adder_tree(2)(425) <= adder_tree(1)(850) + adder_tree(1)(851); --28 bits 
            adder_tree(2)(426) <= adder_tree(1)(852) + adder_tree(1)(853); --28 bits 
            adder_tree(2)(427) <= adder_tree(1)(854) + adder_tree(1)(855); --28 bits 
            adder_tree(2)(428) <= adder_tree(1)(856) + adder_tree(1)(857); --28 bits 
            adder_tree(2)(429) <= adder_tree(1)(858) + adder_tree(1)(859); --28 bits 
            adder_tree(2)(430) <= adder_tree(1)(860) + adder_tree(1)(861); --28 bits 
            adder_tree(2)(431) <= adder_tree(1)(862) + adder_tree(1)(863); --28 bits 
            adder_tree(2)(432) <= adder_tree(1)(864) + adder_tree(1)(865); --28 bits 
            adder_tree(2)(433) <= adder_tree(1)(866) + adder_tree(1)(867); --28 bits 
            adder_tree(2)(434) <= adder_tree(1)(868) + adder_tree(1)(869); --28 bits 
            adder_tree(2)(435) <= adder_tree(1)(870) + adder_tree(1)(871); --28 bits 
            adder_tree(2)(436) <= adder_tree(1)(872) + adder_tree(1)(873); --28 bits 
            adder_tree(2)(437) <= adder_tree(1)(874) + adder_tree(1)(875); --28 bits 
            adder_tree(2)(438) <= adder_tree(1)(876) + adder_tree(1)(877); --28 bits 
            adder_tree(2)(439) <= adder_tree(1)(878) + adder_tree(1)(879); --28 bits 
            adder_tree(2)(440) <= adder_tree(1)(880) + adder_tree(1)(881); --28 bits 
            adder_tree(2)(441) <= adder_tree(1)(882) + adder_tree(1)(883); --28 bits 
            adder_tree(2)(442) <= adder_tree(1)(884) + adder_tree(1)(885); --28 bits 
            adder_tree(2)(443) <= adder_tree(1)(886) + adder_tree(1)(887); --28 bits 
            adder_tree(2)(444) <= adder_tree(1)(888) + adder_tree(1)(889); --28 bits 
            adder_tree(2)(445) <= adder_tree(1)(890) + adder_tree(1)(891); --28 bits 
            adder_tree(2)(446) <= adder_tree(1)(892) + adder_tree(1)(893); --28 bits 
            adder_tree(2)(447) <= adder_tree(1)(894) + adder_tree(1)(895); --28 bits 
            adder_tree(2)(448) <= adder_tree(1)(896) + adder_tree(1)(897); --28 bits 
            adder_tree(2)(449) <= adder_tree(1)(898) + adder_tree(1)(899); --28 bits 
            adder_tree(2)(450) <= adder_tree(1)(900) + adder_tree(1)(901); --28 bits 
            adder_tree(2)(451) <= adder_tree(1)(902) + adder_tree(1)(903); --28 bits 
            adder_tree(2)(452) <= adder_tree(1)(904) + adder_tree(1)(905); --28 bits 
            adder_tree(2)(453) <= adder_tree(1)(906) + adder_tree(1)(907); --28 bits 
            adder_tree(2)(454) <= adder_tree(1)(908) + adder_tree(1)(909); --28 bits 
            adder_tree(2)(455) <= adder_tree(1)(910) + adder_tree(1)(911); --28 bits 
            adder_tree(2)(456) <= adder_tree(1)(912) + adder_tree(1)(913); --28 bits 
            adder_tree(2)(457) <= adder_tree(1)(914) + adder_tree(1)(915); --28 bits 
            adder_tree(2)(458) <= adder_tree(1)(916) + adder_tree(1)(917); --28 bits 
            adder_tree(2)(459) <= adder_tree(1)(918) + adder_tree(1)(919); --28 bits 
            adder_tree(2)(460) <= adder_tree(1)(920) + adder_tree(1)(921); --28 bits 
            adder_tree(2)(461) <= adder_tree(1)(922) + adder_tree(1)(923); --28 bits 
            adder_tree(2)(462) <= adder_tree(1)(924) + adder_tree(1)(925); --28 bits 
            adder_tree(2)(463) <= adder_tree(1)(926) + adder_tree(1)(927); --28 bits 
            adder_tree(2)(464) <= adder_tree(1)(928) + adder_tree(1)(929); --28 bits 
            adder_tree(2)(465) <= adder_tree(1)(930) + adder_tree(1)(931); --28 bits 
            adder_tree(2)(466) <= adder_tree(1)(932) + adder_tree(1)(933); --28 bits 
            adder_tree(2)(467) <= adder_tree(1)(934) + adder_tree(1)(935); --28 bits 
            adder_tree(2)(468) <= adder_tree(1)(936) + adder_tree(1)(937); --28 bits 
            adder_tree(2)(469) <= adder_tree(1)(938) + adder_tree(1)(939); --28 bits 
            adder_tree(2)(470) <= adder_tree(1)(940) + adder_tree(1)(941); --28 bits 
            adder_tree(2)(471) <= adder_tree(1)(942) + adder_tree(1)(943); --28 bits 
            adder_tree(2)(472) <= adder_tree(1)(944) + adder_tree(1)(945); --28 bits 
            adder_tree(2)(473) <= adder_tree(1)(946) + adder_tree(1)(947); --28 bits 
            adder_tree(2)(474) <= adder_tree(1)(948) + adder_tree(1)(949); --28 bits 
            adder_tree(2)(475) <= adder_tree(1)(950) + adder_tree(1)(951); --28 bits 
            adder_tree(2)(476) <= adder_tree(1)(952) + adder_tree(1)(953); --28 bits 
            adder_tree(2)(477) <= adder_tree(1)(954) + adder_tree(1)(955); --28 bits 
            adder_tree(2)(478) <= adder_tree(1)(956) + adder_tree(1)(957); --28 bits 
            adder_tree(2)(479) <= adder_tree(1)(958) + adder_tree(1)(959); --28 bits 
            adder_tree(2)(480) <= adder_tree(1)(960) + adder_tree(1)(961); --28 bits 
            adder_tree(2)(481) <= adder_tree(1)(962) + adder_tree(1)(963); --28 bits 
            adder_tree(2)(482) <= adder_tree(1)(964) + adder_tree(1)(965); --28 bits 
            adder_tree(2)(483) <= adder_tree(1)(966) + adder_tree(1)(967); --28 bits 
            adder_tree(2)(484) <= adder_tree(1)(968) + adder_tree(1)(969); --28 bits 
            adder_tree(2)(485) <= adder_tree(1)(970) + adder_tree(1)(971); --28 bits 
            adder_tree(2)(486) <= adder_tree(1)(972) + adder_tree(1)(973); --28 bits 
            adder_tree(2)(487) <= adder_tree(1)(974) + adder_tree(1)(975); --28 bits 
            adder_tree(2)(488) <= adder_tree(1)(976) + adder_tree(1)(977); --28 bits 
            adder_tree(2)(489) <= adder_tree(1)(978) + adder_tree(1)(979); --28 bits 
            adder_tree(2)(490) <= adder_tree(1)(980) + adder_tree(1)(981); --28 bits 
            adder_tree(2)(491) <= adder_tree(1)(982) + adder_tree(1)(983); --28 bits 
            adder_tree(2)(492) <= adder_tree(1)(984) + adder_tree(1)(985); --28 bits 
            adder_tree(2)(493) <= adder_tree(1)(986) + adder_tree(1)(987); --28 bits 
            adder_tree(2)(494) <= adder_tree(1)(988) + adder_tree(1)(989); --28 bits 
            adder_tree(2)(495) <= adder_tree(1)(990) + adder_tree(1)(991); --28 bits 
            adder_tree(2)(496) <= adder_tree(1)(992) + adder_tree(1)(993); --28 bits 
            adder_tree(2)(497) <= adder_tree(1)(994) + adder_tree(1)(995); --28 bits 
            adder_tree(2)(498) <= adder_tree(1)(996) + adder_tree(1)(997); --28 bits 
            adder_tree(2)(499) <= adder_tree(1)(998) + adder_tree(1)(999); --28 bits 
            adder_tree(2)(500) <= adder_tree(1)(1000) + adder_tree(1)(1001); --28 bits 
            adder_tree(2)(501) <= adder_tree(1)(1002) + adder_tree(1)(1003); --28 bits 
            adder_tree(2)(502) <= adder_tree(1)(1004) + adder_tree(1)(1005); --28 bits 
            adder_tree(2)(503) <= adder_tree(1)(1006) + adder_tree(1)(1007); --28 bits 
            adder_tree(2)(504) <= adder_tree(1)(1008) + adder_tree(1)(1009); --28 bits 
            adder_tree(2)(505) <= adder_tree(1)(1010) + adder_tree(1)(1011); --28 bits 
            adder_tree(2)(506) <= adder_tree(1)(1012) + adder_tree(1)(1013); --28 bits 
            adder_tree(2)(507) <= adder_tree(1)(1014) + adder_tree(1)(1015); --28 bits 
            adder_tree(2)(508) <= adder_tree(1)(1016) + adder_tree(1)(1017); --28 bits 
            adder_tree(2)(509) <= adder_tree(1)(1018) + adder_tree(1)(1019); --28 bits 
            adder_tree(2)(510) <= adder_tree(1)(1020) + adder_tree(1)(1021); --28 bits 
            adder_tree(2)(511) <= adder_tree(1)(1022) + adder_tree(1)(1023); --28 bits 
            adder_tree(2)(512) <= adder_tree(1)(1024) + adder_tree(1)(1025); --28 bits 
            adder_tree(3)(0) <= adder_tree(2)(0) + adder_tree(2)(1); --29 bits 
            adder_tree(3)(1) <= adder_tree(2)(2) + adder_tree(2)(3); --29 bits 
            adder_tree(3)(2) <= adder_tree(2)(4) + adder_tree(2)(5); --29 bits 
            adder_tree(3)(3) <= adder_tree(2)(6) + adder_tree(2)(7); --29 bits 
            adder_tree(3)(4) <= adder_tree(2)(8) + adder_tree(2)(9); --29 bits 
            adder_tree(3)(5) <= adder_tree(2)(10) + adder_tree(2)(11); --29 bits 
            adder_tree(3)(6) <= adder_tree(2)(12) + adder_tree(2)(13); --29 bits 
            adder_tree(3)(7) <= adder_tree(2)(14) + adder_tree(2)(15); --29 bits 
            adder_tree(3)(8) <= adder_tree(2)(16) + adder_tree(2)(17); --29 bits 
            adder_tree(3)(9) <= adder_tree(2)(18) + adder_tree(2)(19); --29 bits 
            adder_tree(3)(10) <= adder_tree(2)(20) + adder_tree(2)(21); --29 bits 
            adder_tree(3)(11) <= adder_tree(2)(22) + adder_tree(2)(23); --29 bits 
            adder_tree(3)(12) <= adder_tree(2)(24) + adder_tree(2)(25); --29 bits 
            adder_tree(3)(13) <= adder_tree(2)(26) + adder_tree(2)(27); --29 bits 
            adder_tree(3)(14) <= adder_tree(2)(28) + adder_tree(2)(29); --29 bits 
            adder_tree(3)(15) <= adder_tree(2)(30) + adder_tree(2)(31); --29 bits 
            adder_tree(3)(16) <= adder_tree(2)(32) + adder_tree(2)(33); --29 bits 
            adder_tree(3)(17) <= adder_tree(2)(34) + adder_tree(2)(35); --29 bits 
            adder_tree(3)(18) <= adder_tree(2)(36) + adder_tree(2)(37); --29 bits 
            adder_tree(3)(19) <= adder_tree(2)(38) + adder_tree(2)(39); --29 bits 
            adder_tree(3)(20) <= adder_tree(2)(40) + adder_tree(2)(41); --29 bits 
            adder_tree(3)(21) <= adder_tree(2)(42) + adder_tree(2)(43); --29 bits 
            adder_tree(3)(22) <= adder_tree(2)(44) + adder_tree(2)(45); --29 bits 
            adder_tree(3)(23) <= adder_tree(2)(46) + adder_tree(2)(47); --29 bits 
            adder_tree(3)(24) <= adder_tree(2)(48) + adder_tree(2)(49); --29 bits 
            adder_tree(3)(25) <= adder_tree(2)(50) + adder_tree(2)(51); --29 bits 
            adder_tree(3)(26) <= adder_tree(2)(52) + adder_tree(2)(53); --29 bits 
            adder_tree(3)(27) <= adder_tree(2)(54) + adder_tree(2)(55); --29 bits 
            adder_tree(3)(28) <= adder_tree(2)(56) + adder_tree(2)(57); --29 bits 
            adder_tree(3)(29) <= adder_tree(2)(58) + adder_tree(2)(59); --29 bits 
            adder_tree(3)(30) <= adder_tree(2)(60) + adder_tree(2)(61); --29 bits 
            adder_tree(3)(31) <= adder_tree(2)(62) + adder_tree(2)(63); --29 bits 
            adder_tree(3)(32) <= adder_tree(2)(64) + adder_tree(2)(65); --29 bits 
            adder_tree(3)(33) <= adder_tree(2)(66) + adder_tree(2)(67); --29 bits 
            adder_tree(3)(34) <= adder_tree(2)(68) + adder_tree(2)(69); --29 bits 
            adder_tree(3)(35) <= adder_tree(2)(70) + adder_tree(2)(71); --29 bits 
            adder_tree(3)(36) <= adder_tree(2)(72) + adder_tree(2)(73); --29 bits 
            adder_tree(3)(37) <= adder_tree(2)(74) + adder_tree(2)(75); --29 bits 
            adder_tree(3)(38) <= adder_tree(2)(76) + adder_tree(2)(77); --29 bits 
            adder_tree(3)(39) <= adder_tree(2)(78) + adder_tree(2)(79); --29 bits 
            adder_tree(3)(40) <= adder_tree(2)(80) + adder_tree(2)(81); --29 bits 
            adder_tree(3)(41) <= adder_tree(2)(82) + adder_tree(2)(83); --29 bits 
            adder_tree(3)(42) <= adder_tree(2)(84) + adder_tree(2)(85); --29 bits 
            adder_tree(3)(43) <= adder_tree(2)(86) + adder_tree(2)(87); --29 bits 
            adder_tree(3)(44) <= adder_tree(2)(88) + adder_tree(2)(89); --29 bits 
            adder_tree(3)(45) <= adder_tree(2)(90) + adder_tree(2)(91); --29 bits 
            adder_tree(3)(46) <= adder_tree(2)(92) + adder_tree(2)(93); --29 bits 
            adder_tree(3)(47) <= adder_tree(2)(94) + adder_tree(2)(95); --29 bits 
            adder_tree(3)(48) <= adder_tree(2)(96) + adder_tree(2)(97); --29 bits 
            adder_tree(3)(49) <= adder_tree(2)(98) + adder_tree(2)(99); --29 bits 
            adder_tree(3)(50) <= adder_tree(2)(100) + adder_tree(2)(101); --29 bits 
            adder_tree(3)(51) <= adder_tree(2)(102) + adder_tree(2)(103); --29 bits 
            adder_tree(3)(52) <= adder_tree(2)(104) + adder_tree(2)(105); --29 bits 
            adder_tree(3)(53) <= adder_tree(2)(106) + adder_tree(2)(107); --29 bits 
            adder_tree(3)(54) <= adder_tree(2)(108) + adder_tree(2)(109); --29 bits 
            adder_tree(3)(55) <= adder_tree(2)(110) + adder_tree(2)(111); --29 bits 
            adder_tree(3)(56) <= adder_tree(2)(112) + adder_tree(2)(113); --29 bits 
            adder_tree(3)(57) <= adder_tree(2)(114) + adder_tree(2)(115); --29 bits 
            adder_tree(3)(58) <= adder_tree(2)(116) + adder_tree(2)(117); --29 bits 
            adder_tree(3)(59) <= adder_tree(2)(118) + adder_tree(2)(119); --29 bits 
            adder_tree(3)(60) <= adder_tree(2)(120) + adder_tree(2)(121); --29 bits 
            adder_tree(3)(61) <= adder_tree(2)(122) + adder_tree(2)(123); --29 bits 
            adder_tree(3)(62) <= adder_tree(2)(124) + adder_tree(2)(125); --29 bits 
            adder_tree(3)(63) <= adder_tree(2)(126) + adder_tree(2)(127); --29 bits 
            adder_tree(3)(64) <= adder_tree(2)(128) + adder_tree(2)(129); --29 bits 
            adder_tree(3)(65) <= adder_tree(2)(130) + adder_tree(2)(131); --29 bits 
            adder_tree(3)(66) <= adder_tree(2)(132) + adder_tree(2)(133); --29 bits 
            adder_tree(3)(67) <= adder_tree(2)(134) + adder_tree(2)(135); --29 bits 
            adder_tree(3)(68) <= adder_tree(2)(136) + adder_tree(2)(137); --29 bits 
            adder_tree(3)(69) <= adder_tree(2)(138) + adder_tree(2)(139); --29 bits 
            adder_tree(3)(70) <= adder_tree(2)(140) + adder_tree(2)(141); --29 bits 
            adder_tree(3)(71) <= adder_tree(2)(142) + adder_tree(2)(143); --29 bits 
            adder_tree(3)(72) <= adder_tree(2)(144) + adder_tree(2)(145); --29 bits 
            adder_tree(3)(73) <= adder_tree(2)(146) + adder_tree(2)(147); --29 bits 
            adder_tree(3)(74) <= adder_tree(2)(148) + adder_tree(2)(149); --29 bits 
            adder_tree(3)(75) <= adder_tree(2)(150) + adder_tree(2)(151); --29 bits 
            adder_tree(3)(76) <= adder_tree(2)(152) + adder_tree(2)(153); --29 bits 
            adder_tree(3)(77) <= adder_tree(2)(154) + adder_tree(2)(155); --29 bits 
            adder_tree(3)(78) <= adder_tree(2)(156) + adder_tree(2)(157); --29 bits 
            adder_tree(3)(79) <= adder_tree(2)(158) + adder_tree(2)(159); --29 bits 
            adder_tree(3)(80) <= adder_tree(2)(160) + adder_tree(2)(161); --29 bits 
            adder_tree(3)(81) <= adder_tree(2)(162) + adder_tree(2)(163); --29 bits 
            adder_tree(3)(82) <= adder_tree(2)(164) + adder_tree(2)(165); --29 bits 
            adder_tree(3)(83) <= adder_tree(2)(166) + adder_tree(2)(167); --29 bits 
            adder_tree(3)(84) <= adder_tree(2)(168) + adder_tree(2)(169); --29 bits 
            adder_tree(3)(85) <= adder_tree(2)(170) + adder_tree(2)(171); --29 bits 
            adder_tree(3)(86) <= adder_tree(2)(172) + adder_tree(2)(173); --29 bits 
            adder_tree(3)(87) <= adder_tree(2)(174) + adder_tree(2)(175); --29 bits 
            adder_tree(3)(88) <= adder_tree(2)(176) + adder_tree(2)(177); --29 bits 
            adder_tree(3)(89) <= adder_tree(2)(178) + adder_tree(2)(179); --29 bits 
            adder_tree(3)(90) <= adder_tree(2)(180) + adder_tree(2)(181); --29 bits 
            adder_tree(3)(91) <= adder_tree(2)(182) + adder_tree(2)(183); --29 bits 
            adder_tree(3)(92) <= adder_tree(2)(184) + adder_tree(2)(185); --29 bits 
            adder_tree(3)(93) <= adder_tree(2)(186) + adder_tree(2)(187); --29 bits 
            adder_tree(3)(94) <= adder_tree(2)(188) + adder_tree(2)(189); --29 bits 
            adder_tree(3)(95) <= adder_tree(2)(190) + adder_tree(2)(191); --29 bits 
            adder_tree(3)(96) <= adder_tree(2)(192) + adder_tree(2)(193); --29 bits 
            adder_tree(3)(97) <= adder_tree(2)(194) + adder_tree(2)(195); --29 bits 
            adder_tree(3)(98) <= adder_tree(2)(196) + adder_tree(2)(197); --29 bits 
            adder_tree(3)(99) <= adder_tree(2)(198) + adder_tree(2)(199); --29 bits 
            adder_tree(3)(100) <= adder_tree(2)(200) + adder_tree(2)(201); --29 bits 
            adder_tree(3)(101) <= adder_tree(2)(202) + adder_tree(2)(203); --29 bits 
            adder_tree(3)(102) <= adder_tree(2)(204) + adder_tree(2)(205); --29 bits 
            adder_tree(3)(103) <= adder_tree(2)(206) + adder_tree(2)(207); --29 bits 
            adder_tree(3)(104) <= adder_tree(2)(208) + adder_tree(2)(209); --29 bits 
            adder_tree(3)(105) <= adder_tree(2)(210) + adder_tree(2)(211); --29 bits 
            adder_tree(3)(106) <= adder_tree(2)(212) + adder_tree(2)(213); --29 bits 
            adder_tree(3)(107) <= adder_tree(2)(214) + adder_tree(2)(215); --29 bits 
            adder_tree(3)(108) <= adder_tree(2)(216) + adder_tree(2)(217); --29 bits 
            adder_tree(3)(109) <= adder_tree(2)(218) + adder_tree(2)(219); --29 bits 
            adder_tree(3)(110) <= adder_tree(2)(220) + adder_tree(2)(221); --29 bits 
            adder_tree(3)(111) <= adder_tree(2)(222) + adder_tree(2)(223); --29 bits 
            adder_tree(3)(112) <= adder_tree(2)(224) + adder_tree(2)(225); --29 bits 
            adder_tree(3)(113) <= adder_tree(2)(226) + adder_tree(2)(227); --29 bits 
            adder_tree(3)(114) <= adder_tree(2)(228) + adder_tree(2)(229); --29 bits 
            adder_tree(3)(115) <= adder_tree(2)(230) + adder_tree(2)(231); --29 bits 
            adder_tree(3)(116) <= adder_tree(2)(232) + adder_tree(2)(233); --29 bits 
            adder_tree(3)(117) <= adder_tree(2)(234) + adder_tree(2)(235); --29 bits 
            adder_tree(3)(118) <= adder_tree(2)(236) + adder_tree(2)(237); --29 bits 
            adder_tree(3)(119) <= adder_tree(2)(238) + adder_tree(2)(239); --29 bits 
            adder_tree(3)(120) <= adder_tree(2)(240) + adder_tree(2)(241); --29 bits 
            adder_tree(3)(121) <= adder_tree(2)(242) + adder_tree(2)(243); --29 bits 
            adder_tree(3)(122) <= adder_tree(2)(244) + adder_tree(2)(245); --29 bits 
            adder_tree(3)(123) <= adder_tree(2)(246) + adder_tree(2)(247); --29 bits 
            adder_tree(3)(124) <= adder_tree(2)(248) + adder_tree(2)(249); --29 bits 
            adder_tree(3)(125) <= adder_tree(2)(250) + adder_tree(2)(251); --29 bits 
            adder_tree(3)(126) <= adder_tree(2)(252) + adder_tree(2)(253); --29 bits 
            adder_tree(3)(127) <= adder_tree(2)(254) + adder_tree(2)(255); --29 bits 
            adder_tree(3)(128) <= adder_tree(2)(256) + adder_tree(2)(257); --29 bits 
            adder_tree(3)(129) <= adder_tree(2)(258) + adder_tree(2)(259); --29 bits 
            adder_tree(3)(130) <= adder_tree(2)(260) + adder_tree(2)(261); --29 bits 
            adder_tree(3)(131) <= adder_tree(2)(262) + adder_tree(2)(263); --29 bits 
            adder_tree(3)(132) <= adder_tree(2)(264) + adder_tree(2)(265); --29 bits 
            adder_tree(3)(133) <= adder_tree(2)(266) + adder_tree(2)(267); --29 bits 
            adder_tree(3)(134) <= adder_tree(2)(268) + adder_tree(2)(269); --29 bits 
            adder_tree(3)(135) <= adder_tree(2)(270) + adder_tree(2)(271); --29 bits 
            adder_tree(3)(136) <= adder_tree(2)(272) + adder_tree(2)(273); --29 bits 
            adder_tree(3)(137) <= adder_tree(2)(274) + adder_tree(2)(275); --29 bits 
            adder_tree(3)(138) <= adder_tree(2)(276) + adder_tree(2)(277); --29 bits 
            adder_tree(3)(139) <= adder_tree(2)(278) + adder_tree(2)(279); --29 bits 
            adder_tree(3)(140) <= adder_tree(2)(280) + adder_tree(2)(281); --29 bits 
            adder_tree(3)(141) <= adder_tree(2)(282) + adder_tree(2)(283); --29 bits 
            adder_tree(3)(142) <= adder_tree(2)(284) + adder_tree(2)(285); --29 bits 
            adder_tree(3)(143) <= adder_tree(2)(286) + adder_tree(2)(287); --29 bits 
            adder_tree(3)(144) <= adder_tree(2)(288) + adder_tree(2)(289); --29 bits 
            adder_tree(3)(145) <= adder_tree(2)(290) + adder_tree(2)(291); --29 bits 
            adder_tree(3)(146) <= adder_tree(2)(292) + adder_tree(2)(293); --29 bits 
            adder_tree(3)(147) <= adder_tree(2)(294) + adder_tree(2)(295); --29 bits 
            adder_tree(3)(148) <= adder_tree(2)(296) + adder_tree(2)(297); --29 bits 
            adder_tree(3)(149) <= adder_tree(2)(298) + adder_tree(2)(299); --29 bits 
            adder_tree(3)(150) <= adder_tree(2)(300) + adder_tree(2)(301); --29 bits 
            adder_tree(3)(151) <= adder_tree(2)(302) + adder_tree(2)(303); --29 bits 
            adder_tree(3)(152) <= adder_tree(2)(304) + adder_tree(2)(305); --29 bits 
            adder_tree(3)(153) <= adder_tree(2)(306) + adder_tree(2)(307); --29 bits 
            adder_tree(3)(154) <= adder_tree(2)(308) + adder_tree(2)(309); --29 bits 
            adder_tree(3)(155) <= adder_tree(2)(310) + adder_tree(2)(311); --29 bits 
            adder_tree(3)(156) <= adder_tree(2)(312) + adder_tree(2)(313); --29 bits 
            adder_tree(3)(157) <= adder_tree(2)(314) + adder_tree(2)(315); --29 bits 
            adder_tree(3)(158) <= adder_tree(2)(316) + adder_tree(2)(317); --29 bits 
            adder_tree(3)(159) <= adder_tree(2)(318) + adder_tree(2)(319); --29 bits 
            adder_tree(3)(160) <= adder_tree(2)(320) + adder_tree(2)(321); --29 bits 
            adder_tree(3)(161) <= adder_tree(2)(322) + adder_tree(2)(323); --29 bits 
            adder_tree(3)(162) <= adder_tree(2)(324) + adder_tree(2)(325); --29 bits 
            adder_tree(3)(163) <= adder_tree(2)(326) + adder_tree(2)(327); --29 bits 
            adder_tree(3)(164) <= adder_tree(2)(328) + adder_tree(2)(329); --29 bits 
            adder_tree(3)(165) <= adder_tree(2)(330) + adder_tree(2)(331); --29 bits 
            adder_tree(3)(166) <= adder_tree(2)(332) + adder_tree(2)(333); --29 bits 
            adder_tree(3)(167) <= adder_tree(2)(334) + adder_tree(2)(335); --29 bits 
            adder_tree(3)(168) <= adder_tree(2)(336) + adder_tree(2)(337); --29 bits 
            adder_tree(3)(169) <= adder_tree(2)(338) + adder_tree(2)(339); --29 bits 
            adder_tree(3)(170) <= adder_tree(2)(340) + adder_tree(2)(341); --29 bits 
            adder_tree(3)(171) <= adder_tree(2)(342) + adder_tree(2)(343); --29 bits 
            adder_tree(3)(172) <= adder_tree(2)(344) + adder_tree(2)(345); --29 bits 
            adder_tree(3)(173) <= adder_tree(2)(346) + adder_tree(2)(347); --29 bits 
            adder_tree(3)(174) <= adder_tree(2)(348) + adder_tree(2)(349); --29 bits 
            adder_tree(3)(175) <= adder_tree(2)(350) + adder_tree(2)(351); --29 bits 
            adder_tree(3)(176) <= adder_tree(2)(352) + adder_tree(2)(353); --29 bits 
            adder_tree(3)(177) <= adder_tree(2)(354) + adder_tree(2)(355); --29 bits 
            adder_tree(3)(178) <= adder_tree(2)(356) + adder_tree(2)(357); --29 bits 
            adder_tree(3)(179) <= adder_tree(2)(358) + adder_tree(2)(359); --29 bits 
            adder_tree(3)(180) <= adder_tree(2)(360) + adder_tree(2)(361); --29 bits 
            adder_tree(3)(181) <= adder_tree(2)(362) + adder_tree(2)(363); --29 bits 
            adder_tree(3)(182) <= adder_tree(2)(364) + adder_tree(2)(365); --29 bits 
            adder_tree(3)(183) <= adder_tree(2)(366) + adder_tree(2)(367); --29 bits 
            adder_tree(3)(184) <= adder_tree(2)(368) + adder_tree(2)(369); --29 bits 
            adder_tree(3)(185) <= adder_tree(2)(370) + adder_tree(2)(371); --29 bits 
            adder_tree(3)(186) <= adder_tree(2)(372) + adder_tree(2)(373); --29 bits 
            adder_tree(3)(187) <= adder_tree(2)(374) + adder_tree(2)(375); --29 bits 
            adder_tree(3)(188) <= adder_tree(2)(376) + adder_tree(2)(377); --29 bits 
            adder_tree(3)(189) <= adder_tree(2)(378) + adder_tree(2)(379); --29 bits 
            adder_tree(3)(190) <= adder_tree(2)(380) + adder_tree(2)(381); --29 bits 
            adder_tree(3)(191) <= adder_tree(2)(382) + adder_tree(2)(383); --29 bits 
            adder_tree(3)(192) <= adder_tree(2)(384) + adder_tree(2)(385); --29 bits 
            adder_tree(3)(193) <= adder_tree(2)(386) + adder_tree(2)(387); --29 bits 
            adder_tree(3)(194) <= adder_tree(2)(388) + adder_tree(2)(389); --29 bits 
            adder_tree(3)(195) <= adder_tree(2)(390) + adder_tree(2)(391); --29 bits 
            adder_tree(3)(196) <= adder_tree(2)(392) + adder_tree(2)(393); --29 bits 
            adder_tree(3)(197) <= adder_tree(2)(394) + adder_tree(2)(395); --29 bits 
            adder_tree(3)(198) <= adder_tree(2)(396) + adder_tree(2)(397); --29 bits 
            adder_tree(3)(199) <= adder_tree(2)(398) + adder_tree(2)(399); --29 bits 
            adder_tree(3)(200) <= adder_tree(2)(400) + adder_tree(2)(401); --29 bits 
            adder_tree(3)(201) <= adder_tree(2)(402) + adder_tree(2)(403); --29 bits 
            adder_tree(3)(202) <= adder_tree(2)(404) + adder_tree(2)(405); --29 bits 
            adder_tree(3)(203) <= adder_tree(2)(406) + adder_tree(2)(407); --29 bits 
            adder_tree(3)(204) <= adder_tree(2)(408) + adder_tree(2)(409); --29 bits 
            adder_tree(3)(205) <= adder_tree(2)(410) + adder_tree(2)(411); --29 bits 
            adder_tree(3)(206) <= adder_tree(2)(412) + adder_tree(2)(413); --29 bits 
            adder_tree(3)(207) <= adder_tree(2)(414) + adder_tree(2)(415); --29 bits 
            adder_tree(3)(208) <= adder_tree(2)(416) + adder_tree(2)(417); --29 bits 
            adder_tree(3)(209) <= adder_tree(2)(418) + adder_tree(2)(419); --29 bits 
            adder_tree(3)(210) <= adder_tree(2)(420) + adder_tree(2)(421); --29 bits 
            adder_tree(3)(211) <= adder_tree(2)(422) + adder_tree(2)(423); --29 bits 
            adder_tree(3)(212) <= adder_tree(2)(424) + adder_tree(2)(425); --29 bits 
            adder_tree(3)(213) <= adder_tree(2)(426) + adder_tree(2)(427); --29 bits 
            adder_tree(3)(214) <= adder_tree(2)(428) + adder_tree(2)(429); --29 bits 
            adder_tree(3)(215) <= adder_tree(2)(430) + adder_tree(2)(431); --29 bits 
            adder_tree(3)(216) <= adder_tree(2)(432) + adder_tree(2)(433); --29 bits 
            adder_tree(3)(217) <= adder_tree(2)(434) + adder_tree(2)(435); --29 bits 
            adder_tree(3)(218) <= adder_tree(2)(436) + adder_tree(2)(437); --29 bits 
            adder_tree(3)(219) <= adder_tree(2)(438) + adder_tree(2)(439); --29 bits 
            adder_tree(3)(220) <= adder_tree(2)(440) + adder_tree(2)(441); --29 bits 
            adder_tree(3)(221) <= adder_tree(2)(442) + adder_tree(2)(443); --29 bits 
            adder_tree(3)(222) <= adder_tree(2)(444) + adder_tree(2)(445); --29 bits 
            adder_tree(3)(223) <= adder_tree(2)(446) + adder_tree(2)(447); --29 bits 
            adder_tree(3)(224) <= adder_tree(2)(448) + adder_tree(2)(449); --29 bits 
            adder_tree(3)(225) <= adder_tree(2)(450) + adder_tree(2)(451); --29 bits 
            adder_tree(3)(226) <= adder_tree(2)(452) + adder_tree(2)(453); --29 bits 
            adder_tree(3)(227) <= adder_tree(2)(454) + adder_tree(2)(455); --29 bits 
            adder_tree(3)(228) <= adder_tree(2)(456) + adder_tree(2)(457); --29 bits 
            adder_tree(3)(229) <= adder_tree(2)(458) + adder_tree(2)(459); --29 bits 
            adder_tree(3)(230) <= adder_tree(2)(460) + adder_tree(2)(461); --29 bits 
            adder_tree(3)(231) <= adder_tree(2)(462) + adder_tree(2)(463); --29 bits 
            adder_tree(3)(232) <= adder_tree(2)(464) + adder_tree(2)(465); --29 bits 
            adder_tree(3)(233) <= adder_tree(2)(466) + adder_tree(2)(467); --29 bits 
            adder_tree(3)(234) <= adder_tree(2)(468) + adder_tree(2)(469); --29 bits 
            adder_tree(3)(235) <= adder_tree(2)(470) + adder_tree(2)(471); --29 bits 
            adder_tree(3)(236) <= adder_tree(2)(472) + adder_tree(2)(473); --29 bits 
            adder_tree(3)(237) <= adder_tree(2)(474) + adder_tree(2)(475); --29 bits 
            adder_tree(3)(238) <= adder_tree(2)(476) + adder_tree(2)(477); --29 bits 
            adder_tree(3)(239) <= adder_tree(2)(478) + adder_tree(2)(479); --29 bits 
            adder_tree(3)(240) <= adder_tree(2)(480) + adder_tree(2)(481); --29 bits 
            adder_tree(3)(241) <= adder_tree(2)(482) + adder_tree(2)(483); --29 bits 
            adder_tree(3)(242) <= adder_tree(2)(484) + adder_tree(2)(485); --29 bits 
            adder_tree(3)(243) <= adder_tree(2)(486) + adder_tree(2)(487); --29 bits 
            adder_tree(3)(244) <= adder_tree(2)(488) + adder_tree(2)(489); --29 bits 
            adder_tree(3)(245) <= adder_tree(2)(490) + adder_tree(2)(491); --29 bits 
            adder_tree(3)(246) <= adder_tree(2)(492) + adder_tree(2)(493); --29 bits 
            adder_tree(3)(247) <= adder_tree(2)(494) + adder_tree(2)(495); --29 bits 
            adder_tree(3)(248) <= adder_tree(2)(496) + adder_tree(2)(497); --29 bits 
            adder_tree(3)(249) <= adder_tree(2)(498) + adder_tree(2)(499); --29 bits 
            adder_tree(3)(250) <= adder_tree(2)(500) + adder_tree(2)(501); --29 bits 
            adder_tree(3)(251) <= adder_tree(2)(502) + adder_tree(2)(503); --29 bits 
            adder_tree(3)(252) <= adder_tree(2)(504) + adder_tree(2)(505); --29 bits 
            adder_tree(3)(253) <= adder_tree(2)(506) + adder_tree(2)(507); --29 bits 
            adder_tree(3)(254) <= adder_tree(2)(508) + adder_tree(2)(509); --29 bits 
            adder_tree(3)(255) <= adder_tree(2)(510) + adder_tree(2)(511); --29 bits 
            adder_tree(3)(256) <= adder_tree(2)(512) + adder_tree(2)(513); --29 bits 
            adder_tree(4)(0) <= adder_tree(3)(0) + adder_tree(3)(1); --30 bits 
            adder_tree(4)(1) <= adder_tree(3)(2) + adder_tree(3)(3); --30 bits 
            adder_tree(4)(2) <= adder_tree(3)(4) + adder_tree(3)(5); --30 bits 
            adder_tree(4)(3) <= adder_tree(3)(6) + adder_tree(3)(7); --30 bits 
            adder_tree(4)(4) <= adder_tree(3)(8) + adder_tree(3)(9); --30 bits 
            adder_tree(4)(5) <= adder_tree(3)(10) + adder_tree(3)(11); --30 bits 
            adder_tree(4)(6) <= adder_tree(3)(12) + adder_tree(3)(13); --30 bits 
            adder_tree(4)(7) <= adder_tree(3)(14) + adder_tree(3)(15); --30 bits 
            adder_tree(4)(8) <= adder_tree(3)(16) + adder_tree(3)(17); --30 bits 
            adder_tree(4)(9) <= adder_tree(3)(18) + adder_tree(3)(19); --30 bits 
            adder_tree(4)(10) <= adder_tree(3)(20) + adder_tree(3)(21); --30 bits 
            adder_tree(4)(11) <= adder_tree(3)(22) + adder_tree(3)(23); --30 bits 
            adder_tree(4)(12) <= adder_tree(3)(24) + adder_tree(3)(25); --30 bits 
            adder_tree(4)(13) <= adder_tree(3)(26) + adder_tree(3)(27); --30 bits 
            adder_tree(4)(14) <= adder_tree(3)(28) + adder_tree(3)(29); --30 bits 
            adder_tree(4)(15) <= adder_tree(3)(30) + adder_tree(3)(31); --30 bits 
            adder_tree(4)(16) <= adder_tree(3)(32) + adder_tree(3)(33); --30 bits 
            adder_tree(4)(17) <= adder_tree(3)(34) + adder_tree(3)(35); --30 bits 
            adder_tree(4)(18) <= adder_tree(3)(36) + adder_tree(3)(37); --30 bits 
            adder_tree(4)(19) <= adder_tree(3)(38) + adder_tree(3)(39); --30 bits 
            adder_tree(4)(20) <= adder_tree(3)(40) + adder_tree(3)(41); --30 bits 
            adder_tree(4)(21) <= adder_tree(3)(42) + adder_tree(3)(43); --30 bits 
            adder_tree(4)(22) <= adder_tree(3)(44) + adder_tree(3)(45); --30 bits 
            adder_tree(4)(23) <= adder_tree(3)(46) + adder_tree(3)(47); --30 bits 
            adder_tree(4)(24) <= adder_tree(3)(48) + adder_tree(3)(49); --30 bits 
            adder_tree(4)(25) <= adder_tree(3)(50) + adder_tree(3)(51); --30 bits 
            adder_tree(4)(26) <= adder_tree(3)(52) + adder_tree(3)(53); --30 bits 
            adder_tree(4)(27) <= adder_tree(3)(54) + adder_tree(3)(55); --30 bits 
            adder_tree(4)(28) <= adder_tree(3)(56) + adder_tree(3)(57); --30 bits 
            adder_tree(4)(29) <= adder_tree(3)(58) + adder_tree(3)(59); --30 bits 
            adder_tree(4)(30) <= adder_tree(3)(60) + adder_tree(3)(61); --30 bits 
            adder_tree(4)(31) <= adder_tree(3)(62) + adder_tree(3)(63); --30 bits 
            adder_tree(4)(32) <= adder_tree(3)(64) + adder_tree(3)(65); --30 bits 
            adder_tree(4)(33) <= adder_tree(3)(66) + adder_tree(3)(67); --30 bits 
            adder_tree(4)(34) <= adder_tree(3)(68) + adder_tree(3)(69); --30 bits 
            adder_tree(4)(35) <= adder_tree(3)(70) + adder_tree(3)(71); --30 bits 
            adder_tree(4)(36) <= adder_tree(3)(72) + adder_tree(3)(73); --30 bits 
            adder_tree(4)(37) <= adder_tree(3)(74) + adder_tree(3)(75); --30 bits 
            adder_tree(4)(38) <= adder_tree(3)(76) + adder_tree(3)(77); --30 bits 
            adder_tree(4)(39) <= adder_tree(3)(78) + adder_tree(3)(79); --30 bits 
            adder_tree(4)(40) <= adder_tree(3)(80) + adder_tree(3)(81); --30 bits 
            adder_tree(4)(41) <= adder_tree(3)(82) + adder_tree(3)(83); --30 bits 
            adder_tree(4)(42) <= adder_tree(3)(84) + adder_tree(3)(85); --30 bits 
            adder_tree(4)(43) <= adder_tree(3)(86) + adder_tree(3)(87); --30 bits 
            adder_tree(4)(44) <= adder_tree(3)(88) + adder_tree(3)(89); --30 bits 
            adder_tree(4)(45) <= adder_tree(3)(90) + adder_tree(3)(91); --30 bits 
            adder_tree(4)(46) <= adder_tree(3)(92) + adder_tree(3)(93); --30 bits 
            adder_tree(4)(47) <= adder_tree(3)(94) + adder_tree(3)(95); --30 bits 
            adder_tree(4)(48) <= adder_tree(3)(96) + adder_tree(3)(97); --30 bits 
            adder_tree(4)(49) <= adder_tree(3)(98) + adder_tree(3)(99); --30 bits 
            adder_tree(4)(50) <= adder_tree(3)(100) + adder_tree(3)(101); --30 bits 
            adder_tree(4)(51) <= adder_tree(3)(102) + adder_tree(3)(103); --30 bits 
            adder_tree(4)(52) <= adder_tree(3)(104) + adder_tree(3)(105); --30 bits 
            adder_tree(4)(53) <= adder_tree(3)(106) + adder_tree(3)(107); --30 bits 
            adder_tree(4)(54) <= adder_tree(3)(108) + adder_tree(3)(109); --30 bits 
            adder_tree(4)(55) <= adder_tree(3)(110) + adder_tree(3)(111); --30 bits 
            adder_tree(4)(56) <= adder_tree(3)(112) + adder_tree(3)(113); --30 bits 
            adder_tree(4)(57) <= adder_tree(3)(114) + adder_tree(3)(115); --30 bits 
            adder_tree(4)(58) <= adder_tree(3)(116) + adder_tree(3)(117); --30 bits 
            adder_tree(4)(59) <= adder_tree(3)(118) + adder_tree(3)(119); --30 bits 
            adder_tree(4)(60) <= adder_tree(3)(120) + adder_tree(3)(121); --30 bits 
            adder_tree(4)(61) <= adder_tree(3)(122) + adder_tree(3)(123); --30 bits 
            adder_tree(4)(62) <= adder_tree(3)(124) + adder_tree(3)(125); --30 bits 
            adder_tree(4)(63) <= adder_tree(3)(126) + adder_tree(3)(127); --30 bits 
            adder_tree(4)(64) <= adder_tree(3)(128) + adder_tree(3)(129); --30 bits 
            adder_tree(4)(65) <= adder_tree(3)(130) + adder_tree(3)(131); --30 bits 
            adder_tree(4)(66) <= adder_tree(3)(132) + adder_tree(3)(133); --30 bits 
            adder_tree(4)(67) <= adder_tree(3)(134) + adder_tree(3)(135); --30 bits 
            adder_tree(4)(68) <= adder_tree(3)(136) + adder_tree(3)(137); --30 bits 
            adder_tree(4)(69) <= adder_tree(3)(138) + adder_tree(3)(139); --30 bits 
            adder_tree(4)(70) <= adder_tree(3)(140) + adder_tree(3)(141); --30 bits 
            adder_tree(4)(71) <= adder_tree(3)(142) + adder_tree(3)(143); --30 bits 
            adder_tree(4)(72) <= adder_tree(3)(144) + adder_tree(3)(145); --30 bits 
            adder_tree(4)(73) <= adder_tree(3)(146) + adder_tree(3)(147); --30 bits 
            adder_tree(4)(74) <= adder_tree(3)(148) + adder_tree(3)(149); --30 bits 
            adder_tree(4)(75) <= adder_tree(3)(150) + adder_tree(3)(151); --30 bits 
            adder_tree(4)(76) <= adder_tree(3)(152) + adder_tree(3)(153); --30 bits 
            adder_tree(4)(77) <= adder_tree(3)(154) + adder_tree(3)(155); --30 bits 
            adder_tree(4)(78) <= adder_tree(3)(156) + adder_tree(3)(157); --30 bits 
            adder_tree(4)(79) <= adder_tree(3)(158) + adder_tree(3)(159); --30 bits 
            adder_tree(4)(80) <= adder_tree(3)(160) + adder_tree(3)(161); --30 bits 
            adder_tree(4)(81) <= adder_tree(3)(162) + adder_tree(3)(163); --30 bits 
            adder_tree(4)(82) <= adder_tree(3)(164) + adder_tree(3)(165); --30 bits 
            adder_tree(4)(83) <= adder_tree(3)(166) + adder_tree(3)(167); --30 bits 
            adder_tree(4)(84) <= adder_tree(3)(168) + adder_tree(3)(169); --30 bits 
            adder_tree(4)(85) <= adder_tree(3)(170) + adder_tree(3)(171); --30 bits 
            adder_tree(4)(86) <= adder_tree(3)(172) + adder_tree(3)(173); --30 bits 
            adder_tree(4)(87) <= adder_tree(3)(174) + adder_tree(3)(175); --30 bits 
            adder_tree(4)(88) <= adder_tree(3)(176) + adder_tree(3)(177); --30 bits 
            adder_tree(4)(89) <= adder_tree(3)(178) + adder_tree(3)(179); --30 bits 
            adder_tree(4)(90) <= adder_tree(3)(180) + adder_tree(3)(181); --30 bits 
            adder_tree(4)(91) <= adder_tree(3)(182) + adder_tree(3)(183); --30 bits 
            adder_tree(4)(92) <= adder_tree(3)(184) + adder_tree(3)(185); --30 bits 
            adder_tree(4)(93) <= adder_tree(3)(186) + adder_tree(3)(187); --30 bits 
            adder_tree(4)(94) <= adder_tree(3)(188) + adder_tree(3)(189); --30 bits 
            adder_tree(4)(95) <= adder_tree(3)(190) + adder_tree(3)(191); --30 bits 
            adder_tree(4)(96) <= adder_tree(3)(192) + adder_tree(3)(193); --30 bits 
            adder_tree(4)(97) <= adder_tree(3)(194) + adder_tree(3)(195); --30 bits 
            adder_tree(4)(98) <= adder_tree(3)(196) + adder_tree(3)(197); --30 bits 
            adder_tree(4)(99) <= adder_tree(3)(198) + adder_tree(3)(199); --30 bits 
            adder_tree(4)(100) <= adder_tree(3)(200) + adder_tree(3)(201); --30 bits 
            adder_tree(4)(101) <= adder_tree(3)(202) + adder_tree(3)(203); --30 bits 
            adder_tree(4)(102) <= adder_tree(3)(204) + adder_tree(3)(205); --30 bits 
            adder_tree(4)(103) <= adder_tree(3)(206) + adder_tree(3)(207); --30 bits 
            adder_tree(4)(104) <= adder_tree(3)(208) + adder_tree(3)(209); --30 bits 
            adder_tree(4)(105) <= adder_tree(3)(210) + adder_tree(3)(211); --30 bits 
            adder_tree(4)(106) <= adder_tree(3)(212) + adder_tree(3)(213); --30 bits 
            adder_tree(4)(107) <= adder_tree(3)(214) + adder_tree(3)(215); --30 bits 
            adder_tree(4)(108) <= adder_tree(3)(216) + adder_tree(3)(217); --30 bits 
            adder_tree(4)(109) <= adder_tree(3)(218) + adder_tree(3)(219); --30 bits 
            adder_tree(4)(110) <= adder_tree(3)(220) + adder_tree(3)(221); --30 bits 
            adder_tree(4)(111) <= adder_tree(3)(222) + adder_tree(3)(223); --30 bits 
            adder_tree(4)(112) <= adder_tree(3)(224) + adder_tree(3)(225); --30 bits 
            adder_tree(4)(113) <= adder_tree(3)(226) + adder_tree(3)(227); --30 bits 
            adder_tree(4)(114) <= adder_tree(3)(228) + adder_tree(3)(229); --30 bits 
            adder_tree(4)(115) <= adder_tree(3)(230) + adder_tree(3)(231); --30 bits 
            adder_tree(4)(116) <= adder_tree(3)(232) + adder_tree(3)(233); --30 bits 
            adder_tree(4)(117) <= adder_tree(3)(234) + adder_tree(3)(235); --30 bits 
            adder_tree(4)(118) <= adder_tree(3)(236) + adder_tree(3)(237); --30 bits 
            adder_tree(4)(119) <= adder_tree(3)(238) + adder_tree(3)(239); --30 bits 
            adder_tree(4)(120) <= adder_tree(3)(240) + adder_tree(3)(241); --30 bits 
            adder_tree(4)(121) <= adder_tree(3)(242) + adder_tree(3)(243); --30 bits 
            adder_tree(4)(122) <= adder_tree(3)(244) + adder_tree(3)(245); --30 bits 
            adder_tree(4)(123) <= adder_tree(3)(246) + adder_tree(3)(247); --30 bits 
            adder_tree(4)(124) <= adder_tree(3)(248) + adder_tree(3)(249); --30 bits 
            adder_tree(4)(125) <= adder_tree(3)(250) + adder_tree(3)(251); --30 bits 
            adder_tree(4)(126) <= adder_tree(3)(252) + adder_tree(3)(253); --30 bits 
            adder_tree(4)(127) <= adder_tree(3)(254) + adder_tree(3)(255); --30 bits 
            adder_tree(4)(128) <= adder_tree(3)(256) + adder_tree(3)(257); --30 bits 
            adder_tree(5)(0) <= adder_tree(4)(0) + adder_tree(4)(1); --31 bits 
            adder_tree(5)(1) <= adder_tree(4)(2) + adder_tree(4)(3); --31 bits 
            adder_tree(5)(2) <= adder_tree(4)(4) + adder_tree(4)(5); --31 bits 
            adder_tree(5)(3) <= adder_tree(4)(6) + adder_tree(4)(7); --31 bits 
            adder_tree(5)(4) <= adder_tree(4)(8) + adder_tree(4)(9); --31 bits 
            adder_tree(5)(5) <= adder_tree(4)(10) + adder_tree(4)(11); --31 bits 
            adder_tree(5)(6) <= adder_tree(4)(12) + adder_tree(4)(13); --31 bits 
            adder_tree(5)(7) <= adder_tree(4)(14) + adder_tree(4)(15); --31 bits 
            adder_tree(5)(8) <= adder_tree(4)(16) + adder_tree(4)(17); --31 bits 
            adder_tree(5)(9) <= adder_tree(4)(18) + adder_tree(4)(19); --31 bits 
            adder_tree(5)(10) <= adder_tree(4)(20) + adder_tree(4)(21); --31 bits 
            adder_tree(5)(11) <= adder_tree(4)(22) + adder_tree(4)(23); --31 bits 
            adder_tree(5)(12) <= adder_tree(4)(24) + adder_tree(4)(25); --31 bits 
            adder_tree(5)(13) <= adder_tree(4)(26) + adder_tree(4)(27); --31 bits 
            adder_tree(5)(14) <= adder_tree(4)(28) + adder_tree(4)(29); --31 bits 
            adder_tree(5)(15) <= adder_tree(4)(30) + adder_tree(4)(31); --31 bits 
            adder_tree(5)(16) <= adder_tree(4)(32) + adder_tree(4)(33); --31 bits 
            adder_tree(5)(17) <= adder_tree(4)(34) + adder_tree(4)(35); --31 bits 
            adder_tree(5)(18) <= adder_tree(4)(36) + adder_tree(4)(37); --31 bits 
            adder_tree(5)(19) <= adder_tree(4)(38) + adder_tree(4)(39); --31 bits 
            adder_tree(5)(20) <= adder_tree(4)(40) + adder_tree(4)(41); --31 bits 
            adder_tree(5)(21) <= adder_tree(4)(42) + adder_tree(4)(43); --31 bits 
            adder_tree(5)(22) <= adder_tree(4)(44) + adder_tree(4)(45); --31 bits 
            adder_tree(5)(23) <= adder_tree(4)(46) + adder_tree(4)(47); --31 bits 
            adder_tree(5)(24) <= adder_tree(4)(48) + adder_tree(4)(49); --31 bits 
            adder_tree(5)(25) <= adder_tree(4)(50) + adder_tree(4)(51); --31 bits 
            adder_tree(5)(26) <= adder_tree(4)(52) + adder_tree(4)(53); --31 bits 
            adder_tree(5)(27) <= adder_tree(4)(54) + adder_tree(4)(55); --31 bits 
            adder_tree(5)(28) <= adder_tree(4)(56) + adder_tree(4)(57); --31 bits 
            adder_tree(5)(29) <= adder_tree(4)(58) + adder_tree(4)(59); --31 bits 
            adder_tree(5)(30) <= adder_tree(4)(60) + adder_tree(4)(61); --31 bits 
            adder_tree(5)(31) <= adder_tree(4)(62) + adder_tree(4)(63); --31 bits 
            adder_tree(5)(32) <= adder_tree(4)(64) + adder_tree(4)(65); --31 bits 
            adder_tree(5)(33) <= adder_tree(4)(66) + adder_tree(4)(67); --31 bits 
            adder_tree(5)(34) <= adder_tree(4)(68) + adder_tree(4)(69); --31 bits 
            adder_tree(5)(35) <= adder_tree(4)(70) + adder_tree(4)(71); --31 bits 
            adder_tree(5)(36) <= adder_tree(4)(72) + adder_tree(4)(73); --31 bits 
            adder_tree(5)(37) <= adder_tree(4)(74) + adder_tree(4)(75); --31 bits 
            adder_tree(5)(38) <= adder_tree(4)(76) + adder_tree(4)(77); --31 bits 
            adder_tree(5)(39) <= adder_tree(4)(78) + adder_tree(4)(79); --31 bits 
            adder_tree(5)(40) <= adder_tree(4)(80) + adder_tree(4)(81); --31 bits 
            adder_tree(5)(41) <= adder_tree(4)(82) + adder_tree(4)(83); --31 bits 
            adder_tree(5)(42) <= adder_tree(4)(84) + adder_tree(4)(85); --31 bits 
            adder_tree(5)(43) <= adder_tree(4)(86) + adder_tree(4)(87); --31 bits 
            adder_tree(5)(44) <= adder_tree(4)(88) + adder_tree(4)(89); --31 bits 
            adder_tree(5)(45) <= adder_tree(4)(90) + adder_tree(4)(91); --31 bits 
            adder_tree(5)(46) <= adder_tree(4)(92) + adder_tree(4)(93); --31 bits 
            adder_tree(5)(47) <= adder_tree(4)(94) + adder_tree(4)(95); --31 bits 
            adder_tree(5)(48) <= adder_tree(4)(96) + adder_tree(4)(97); --31 bits 
            adder_tree(5)(49) <= adder_tree(4)(98) + adder_tree(4)(99); --31 bits 
            adder_tree(5)(50) <= adder_tree(4)(100) + adder_tree(4)(101); --31 bits 
            adder_tree(5)(51) <= adder_tree(4)(102) + adder_tree(4)(103); --31 bits 
            adder_tree(5)(52) <= adder_tree(4)(104) + adder_tree(4)(105); --31 bits 
            adder_tree(5)(53) <= adder_tree(4)(106) + adder_tree(4)(107); --31 bits 
            adder_tree(5)(54) <= adder_tree(4)(108) + adder_tree(4)(109); --31 bits 
            adder_tree(5)(55) <= adder_tree(4)(110) + adder_tree(4)(111); --31 bits 
            adder_tree(5)(56) <= adder_tree(4)(112) + adder_tree(4)(113); --31 bits 
            adder_tree(5)(57) <= adder_tree(4)(114) + adder_tree(4)(115); --31 bits 
            adder_tree(5)(58) <= adder_tree(4)(116) + adder_tree(4)(117); --31 bits 
            adder_tree(5)(59) <= adder_tree(4)(118) + adder_tree(4)(119); --31 bits 
            adder_tree(5)(60) <= adder_tree(4)(120) + adder_tree(4)(121); --31 bits 
            adder_tree(5)(61) <= adder_tree(4)(122) + adder_tree(4)(123); --31 bits 
            adder_tree(5)(62) <= adder_tree(4)(124) + adder_tree(4)(125); --31 bits 
            adder_tree(5)(63) <= adder_tree(4)(126) + adder_tree(4)(127); --31 bits 
            adder_tree(5)(64) <= adder_tree(4)(128) + adder_tree(4)(129); --31 bits 
            adder_tree(6)(0) <= adder_tree(5)(0) + adder_tree(5)(1); --32 bits 
            adder_tree(6)(1) <= adder_tree(5)(2) + adder_tree(5)(3); --32 bits 
            adder_tree(6)(2) <= adder_tree(5)(4) + adder_tree(5)(5); --32 bits 
            adder_tree(6)(3) <= adder_tree(5)(6) + adder_tree(5)(7); --32 bits 
            adder_tree(6)(4) <= adder_tree(5)(8) + adder_tree(5)(9); --32 bits 
            adder_tree(6)(5) <= adder_tree(5)(10) + adder_tree(5)(11); --32 bits 
            adder_tree(6)(6) <= adder_tree(5)(12) + adder_tree(5)(13); --32 bits 
            adder_tree(6)(7) <= adder_tree(5)(14) + adder_tree(5)(15); --32 bits 
            adder_tree(6)(8) <= adder_tree(5)(16) + adder_tree(5)(17); --32 bits 
            adder_tree(6)(9) <= adder_tree(5)(18) + adder_tree(5)(19); --32 bits 
            adder_tree(6)(10) <= adder_tree(5)(20) + adder_tree(5)(21); --32 bits 
            adder_tree(6)(11) <= adder_tree(5)(22) + adder_tree(5)(23); --32 bits 
            adder_tree(6)(12) <= adder_tree(5)(24) + adder_tree(5)(25); --32 bits 
            adder_tree(6)(13) <= adder_tree(5)(26) + adder_tree(5)(27); --32 bits 
            adder_tree(6)(14) <= adder_tree(5)(28) + adder_tree(5)(29); --32 bits 
            adder_tree(6)(15) <= adder_tree(5)(30) + adder_tree(5)(31); --32 bits 
            adder_tree(6)(16) <= adder_tree(5)(32) + adder_tree(5)(33); --32 bits 
            adder_tree(6)(17) <= adder_tree(5)(34) + adder_tree(5)(35); --32 bits 
            adder_tree(6)(18) <= adder_tree(5)(36) + adder_tree(5)(37); --32 bits 
            adder_tree(6)(19) <= adder_tree(5)(38) + adder_tree(5)(39); --32 bits 
            adder_tree(6)(20) <= adder_tree(5)(40) + adder_tree(5)(41); --32 bits 
            adder_tree(6)(21) <= adder_tree(5)(42) + adder_tree(5)(43); --32 bits 
            adder_tree(6)(22) <= adder_tree(5)(44) + adder_tree(5)(45); --32 bits 
            adder_tree(6)(23) <= adder_tree(5)(46) + adder_tree(5)(47); --32 bits 
            adder_tree(6)(24) <= adder_tree(5)(48) + adder_tree(5)(49); --32 bits 
            adder_tree(6)(25) <= adder_tree(5)(50) + adder_tree(5)(51); --32 bits 
            adder_tree(6)(26) <= adder_tree(5)(52) + adder_tree(5)(53); --32 bits 
            adder_tree(6)(27) <= adder_tree(5)(54) + adder_tree(5)(55); --32 bits 
            adder_tree(6)(28) <= adder_tree(5)(56) + adder_tree(5)(57); --32 bits 
            adder_tree(6)(29) <= adder_tree(5)(58) + adder_tree(5)(59); --32 bits 
            adder_tree(6)(30) <= adder_tree(5)(60) + adder_tree(5)(61); --32 bits 
            adder_tree(6)(31) <= adder_tree(5)(62) + adder_tree(5)(63); --32 bits 
            adder_tree(6)(32) <= adder_tree(5)(64) + adder_tree(5)(65); --32 bits 
            adder_tree(7)(0) <= adder_tree(6)(0) + adder_tree(6)(1); --33 bits 
            adder_tree(7)(1) <= adder_tree(6)(2) + adder_tree(6)(3); --33 bits 
            adder_tree(7)(2) <= adder_tree(6)(4) + adder_tree(6)(5); --33 bits 
            adder_tree(7)(3) <= adder_tree(6)(6) + adder_tree(6)(7); --33 bits 
            adder_tree(7)(4) <= adder_tree(6)(8) + adder_tree(6)(9); --33 bits 
            adder_tree(7)(5) <= adder_tree(6)(10) + adder_tree(6)(11); --33 bits 
            adder_tree(7)(6) <= adder_tree(6)(12) + adder_tree(6)(13); --33 bits 
            adder_tree(7)(7) <= adder_tree(6)(14) + adder_tree(6)(15); --33 bits 
            adder_tree(7)(8) <= adder_tree(6)(16) + adder_tree(6)(17); --33 bits 
            adder_tree(7)(9) <= adder_tree(6)(18) + adder_tree(6)(19); --33 bits 
            adder_tree(7)(10) <= adder_tree(6)(20) + adder_tree(6)(21); --33 bits 
            adder_tree(7)(11) <= adder_tree(6)(22) + adder_tree(6)(23); --33 bits 
            adder_tree(7)(12) <= adder_tree(6)(24) + adder_tree(6)(25); --33 bits 
            adder_tree(7)(13) <= adder_tree(6)(26) + adder_tree(6)(27); --33 bits 
            adder_tree(7)(14) <= adder_tree(6)(28) + adder_tree(6)(29); --33 bits 
            adder_tree(7)(15) <= adder_tree(6)(30) + adder_tree(6)(31); --33 bits 
            adder_tree(7)(16) <= adder_tree(6)(32) + adder_tree(6)(33); --33 bits 
            adder_tree(8)(0) <= adder_tree(7)(0) + adder_tree(7)(1); --34 bits 
            adder_tree(8)(1) <= adder_tree(7)(2) + adder_tree(7)(3); --34 bits 
            adder_tree(8)(2) <= adder_tree(7)(4) + adder_tree(7)(5); --34 bits 
            adder_tree(8)(3) <= adder_tree(7)(6) + adder_tree(7)(7); --34 bits 
            adder_tree(8)(4) <= adder_tree(7)(8) + adder_tree(7)(9); --34 bits 
            adder_tree(8)(5) <= adder_tree(7)(10) + adder_tree(7)(11); --34 bits 
            adder_tree(8)(6) <= adder_tree(7)(12) + adder_tree(7)(13); --34 bits 
            adder_tree(8)(7) <= adder_tree(7)(14) + adder_tree(7)(15); --34 bits 
            adder_tree(8)(8) <= adder_tree(7)(16) + adder_tree(7)(17); --34 bits 
            adder_tree(9)(0) <= adder_tree(8)(0) + adder_tree(8)(1); --35 bits 
            adder_tree(9)(1) <= adder_tree(8)(2) + adder_tree(8)(3); --35 bits 
            adder_tree(9)(2) <= adder_tree(8)(4) + adder_tree(8)(5); --35 bits 
            adder_tree(9)(3) <= adder_tree(8)(6) + adder_tree(8)(7); --35 bits 
            adder_tree(9)(4) <= adder_tree(8)(8) + adder_tree(8)(9); --35 bits 
            adder_tree(10)(0) <= adder_tree(9)(0) + adder_tree(9)(1); --36 bits 
            adder_tree(10)(1) <= adder_tree(9)(2) + adder_tree(9)(3); --36 bits 
            adder_tree(10)(2) <= adder_tree(9)(4) + adder_tree(9)(5); --36 bits 
            adder_tree(11)(0) <= adder_tree(10)(0) + adder_tree(10)(1);
                                                                                                         
            v_round := '0' & adder_tree(11)(0)(15.0001);                                                     
            data_out_prepare <= std_logic_vector(adder_tree(11)(0)(27.0001 downto 16.0001) + v_round);                                                                         
            data_out_prepare_en <= adder_tree_en(11);                                                    
                                                                                                         
                                                                                                         
                                                                                                         
            adder_tree_en(0) <= data_in_en_r2;                                                           
            adder_tree_en(nb_taps-1 downto 1) <= adder_tree_en(nb_taps-2 downto 0);                      
                                                                                                         
       end if;                                                                                           
    end process;                                                                                         
                                                                                                         
                                                                                                         
                                                                                                         
 data_out     <= data_out_prepare;                                                                       
 data_out_en  <= data_out_prepare_en;                                                                    
                                                                                                         
                                                                                                         
                                                                                                         
 taps(0) <= to_signed(0,14);
 taps(1) <= to_signed(0,14);
 taps(2) <= to_signed(0,14);
 taps(3) <= to_signed(0,14);
 taps(4) <= to_signed(0,14);
 taps(5) <= to_signed(0,14);
 taps(6) <= to_signed(0,14);
 taps(7) <= to_signed(0,14);
 taps(8) <= to_signed(0,14);
 taps(9) <= to_signed(0,14);
 taps(10) <= to_signed(0,14);
 taps(11) <= to_signed(0,14);
 taps(12) <= to_signed(0,14);
 taps(13) <= to_signed(0,14);
 taps(14) <= to_signed(0,14);
 taps(15) <= to_signed(0,14);
 taps(16) <= to_signed(0,14);
 taps(17) <= to_signed(0,14);
 taps(18) <= to_signed(0,14);
 taps(19) <= to_signed(0,14);
 taps(20) <= to_signed(0,14);
 taps(21) <= to_signed(0,14);
 taps(22) <= to_signed(0,14);
 taps(23) <= to_signed(0,14);
 taps(24) <= to_signed(0,14);
 taps(25) <= to_signed(0,14);
 taps(26) <= to_signed(0,14);
 taps(27) <= to_signed(0,14);
 taps(28) <= to_signed(0,14);
 taps(29) <= to_signed(0,14);
 taps(30) <= to_signed(0,14);
 taps(31) <= to_signed(0,14);
 taps(32) <= to_signed(0,14);
 taps(33) <= to_signed(0,14);
 taps(34) <= to_signed(0,14);
 taps(35) <= to_signed(0,14);
 taps(36) <= to_signed(0,14);
 taps(37) <= to_signed(0,14);
 taps(38) <= to_signed(0,14);
 taps(39) <= to_signed(0,14);
 taps(40) <= to_signed(0,14);
 taps(41) <= to_signed(0,14);
 taps(42) <= to_signed(0,14);
 taps(43) <= to_signed(0,14);
 taps(44) <= to_signed(0,14);
 taps(45) <= to_signed(0,14);
 taps(46) <= to_signed(0,14);
 taps(47) <= to_signed(0,14);
 taps(48) <= to_signed(0,14);
 taps(49) <= to_signed(0,14);
 taps(50) <= to_signed(0,14);
 taps(51) <= to_signed(0,14);
 taps(52) <= to_signed(0,14);
 taps(53) <= to_signed(0,14);
 taps(54) <= to_signed(0,14);
 taps(55) <= to_signed(0,14);
 taps(56) <= to_signed(0,14);
 taps(57) <= to_signed(0,14);
 taps(58) <= to_signed(0,14);
 taps(59) <= to_signed(0,14);
 taps(60) <= to_signed(0,14);
 taps(61) <= to_signed(0,14);
 taps(62) <= to_signed(0,14);
 taps(63) <= to_signed(0,14);
 taps(64) <= to_signed(0,14);
 taps(65) <= to_signed(0,14);
 taps(66) <= to_signed(0,14);
 taps(67) <= to_signed(0,14);
 taps(68) <= to_signed(0,14);
 taps(69) <= to_signed(0,14);
 taps(70) <= to_signed(0,14);
 taps(71) <= to_signed(0,14);
 taps(72) <= to_signed(0,14);
 taps(73) <= to_signed(0,14);
 taps(74) <= to_signed(0,14);
 taps(75) <= to_signed(0,14);
 taps(76) <= to_signed(0,14);
 taps(77) <= to_signed(0,14);
 taps(78) <= to_signed(0,14);
 taps(79) <= to_signed(0,14);
 taps(80) <= to_signed(0,14);
 taps(81) <= to_signed(0,14);
 taps(82) <= to_signed(0,14);
 taps(83) <= to_signed(0,14);
 taps(84) <= to_signed(0,14);
 taps(85) <= to_signed(0,14);
 taps(86) <= to_signed(0,14);
 taps(87) <= to_signed(0,14);
 taps(88) <= to_signed(0,14);
 taps(89) <= to_signed(0,14);
 taps(90) <= to_signed(0,14);
 taps(91) <= to_signed(0,14);
 taps(92) <= to_signed(0,14);
 taps(93) <= to_signed(0,14);
 taps(94) <= to_signed(0,14);
 taps(95) <= to_signed(0,14);
 taps(96) <= to_signed(0,14);
 taps(97) <= to_signed(0,14);
 taps(98) <= to_signed(0,14);
 taps(99) <= to_signed(0,14);
 taps(100) <= to_signed(0,14);
 taps(101) <= to_signed(0,14);
 taps(102) <= to_signed(0,14);
 taps(103) <= to_signed(0,14);
 taps(104) <= to_signed(0,14);
 taps(105) <= to_signed(0,14);
 taps(106) <= to_signed(0,14);
 taps(107) <= to_signed(0,14);
 taps(108) <= to_signed(0,14);
 taps(109) <= to_signed(0,14);
 taps(110) <= to_signed(0,14);
 taps(111) <= to_signed(0,14);
 taps(112) <= to_signed(0,14);
 taps(113) <= to_signed(0,14);
 taps(114) <= to_signed(0,14);
 taps(115) <= to_signed(0,14);
 taps(116) <= to_signed(0,14);
 taps(117) <= to_signed(0,14);
 taps(118) <= to_signed(0,14);
 taps(119) <= to_signed(0,14);
 taps(120) <= to_signed(0,14);
 taps(121) <= to_signed(0,14);
 taps(122) <= to_signed(0,14);
 taps(123) <= to_signed(0,14);
 taps(124) <= to_signed(0,14);
 taps(125) <= to_signed(0,14);
 taps(126) <= to_signed(0,14);
 taps(127) <= to_signed(0,14);
 taps(128) <= to_signed(0,14);
 taps(129) <= to_signed(0,14);
 taps(130) <= to_signed(0,14);
 taps(131) <= to_signed(0,14);
 taps(132) <= to_signed(0,14);
 taps(133) <= to_signed(0,14);
 taps(134) <= to_signed(0,14);
 taps(135) <= to_signed(0,14);
 taps(136) <= to_signed(0,14);
 taps(137) <= to_signed(0,14);
 taps(138) <= to_signed(0,14);
 taps(139) <= to_signed(0,14);
 taps(140) <= to_signed(0,14);
 taps(141) <= to_signed(0,14);
 taps(142) <= to_signed(0,14);
 taps(143) <= to_signed(0,14);
 taps(144) <= to_signed(0,14);
 taps(145) <= to_signed(0,14);
 taps(146) <= to_signed(0,14);
 taps(147) <= to_signed(0,14);
 taps(148) <= to_signed(0,14);
 taps(149) <= to_signed(0,14);
 taps(150) <= to_signed(0,14);
 taps(151) <= to_signed(0,14);
 taps(152) <= to_signed(0,14);
 taps(153) <= to_signed(0,14);
 taps(154) <= to_signed(0,14);
 taps(155) <= to_signed(0,14);
 taps(156) <= to_signed(0,14);
 taps(157) <= to_signed(0,14);
 taps(158) <= to_signed(0,14);
 taps(159) <= to_signed(0,14);
 taps(160) <= to_signed(0,14);
 taps(161) <= to_signed(0,14);
 taps(162) <= to_signed(0,14);
 taps(163) <= to_signed(0,14);
 taps(164) <= to_signed(0,14);
 taps(165) <= to_signed(0,14);
 taps(166) <= to_signed(0,14);
 taps(167) <= to_signed(0,14);
 taps(168) <= to_signed(0,14);
 taps(169) <= to_signed(0,14);
 taps(170) <= to_signed(0,14);
 taps(171) <= to_signed(0,14);
 taps(172) <= to_signed(0,14);
 taps(173) <= to_signed(0,14);
 taps(174) <= to_signed(0,14);
 taps(175) <= to_signed(0,14);
 taps(176) <= to_signed(0,14);
 taps(177) <= to_signed(0,14);
 taps(178) <= to_signed(0,14);
 taps(179) <= to_signed(0,14);
 taps(180) <= to_signed(0,14);
 taps(181) <= to_signed(0,14);
 taps(182) <= to_signed(0,14);
 taps(183) <= to_signed(0,14);
 taps(184) <= to_signed(0,14);
 taps(185) <= to_signed(0,14);
 taps(186) <= to_signed(0,14);
 taps(187) <= to_signed(0,14);
 taps(188) <= to_signed(0,14);
 taps(189) <= to_signed(0,14);
 taps(190) <= to_signed(0,14);
 taps(191) <= to_signed(0,14);
 taps(192) <= to_signed(0,14);
 taps(193) <= to_signed(0,14);
 taps(194) <= to_signed(0,14);
 taps(195) <= to_signed(0,14);
 taps(196) <= to_signed(0,14);
 taps(197) <= to_signed(0,14);
 taps(198) <= to_signed(0,14);
 taps(199) <= to_signed(0,14);
 taps(200) <= to_signed(0,14);
 taps(201) <= to_signed(0,14);
 taps(202) <= to_signed(0,14);
 taps(203) <= to_signed(0,14);
 taps(204) <= to_signed(0,14);
 taps(205) <= to_signed(0,14);
 taps(206) <= to_signed(0,14);
 taps(207) <= to_signed(0,14);
 taps(208) <= to_signed(0,14);
 taps(209) <= to_signed(0,14);
 taps(210) <= to_signed(0,14);
 taps(211) <= to_signed(0,14);
 taps(212) <= to_signed(0,14);
 taps(213) <= to_signed(0,14);
 taps(214) <= to_signed(0,14);
 taps(215) <= to_signed(0,14);
 taps(216) <= to_signed(0,14);
 taps(217) <= to_signed(0,14);
 taps(218) <= to_signed(0,14);
 taps(219) <= to_signed(0,14);
 taps(220) <= to_signed(0,14);
 taps(221) <= to_signed(0,14);
 taps(222) <= to_signed(0,14);
 taps(223) <= to_signed(0,14);
 taps(224) <= to_signed(0,14);
 taps(225) <= to_signed(0,14);
 taps(226) <= to_signed(0,14);
 taps(227) <= to_signed(0,14);
 taps(228) <= to_signed(0,14);
 taps(229) <= to_signed(0,14);
 taps(230) <= to_signed(0,14);
 taps(231) <= to_signed(0,14);
 taps(232) <= to_signed(0,14);
 taps(233) <= to_signed(0,14);
 taps(234) <= to_signed(0,14);
 taps(235) <= to_signed(0,14);
 taps(236) <= to_signed(0,14);
 taps(237) <= to_signed(0,14);
 taps(238) <= to_signed(0,14);
 taps(239) <= to_signed(0,14);
 taps(240) <= to_signed(0,14);
 taps(241) <= to_signed(0,14);
 taps(242) <= to_signed(0,14);
 taps(243) <= to_signed(0,14);
 taps(244) <= to_signed(0,14);
 taps(245) <= to_signed(0,14);
 taps(246) <= to_signed(0,14);
 taps(247) <= to_signed(0,14);
 taps(248) <= to_signed(0,14);
 taps(249) <= to_signed(0,14);
 taps(250) <= to_signed(0,14);
 taps(251) <= to_signed(0,14);
 taps(252) <= to_signed(0,14);
 taps(253) <= to_signed(0,14);
 taps(254) <= to_signed(0,14);
 taps(255) <= to_signed(0,14);
 taps(256) <= to_signed(0,14);
 taps(257) <= to_signed(0,14);
 taps(258) <= to_signed(0,14);
 taps(259) <= to_signed(0,14);
 taps(260) <= to_signed(0,14);
 taps(261) <= to_signed(0,14);
 taps(262) <= to_signed(0,14);
 taps(263) <= to_signed(0,14);
 taps(264) <= to_signed(0,14);
 taps(265) <= to_signed(0,14);
 taps(266) <= to_signed(0,14);
 taps(267) <= to_signed(0,14);
 taps(268) <= to_signed(0,14);
 taps(269) <= to_signed(0,14);
 taps(270) <= to_signed(0,14);
 taps(271) <= to_signed(0,14);
 taps(272) <= to_signed(0,14);
 taps(273) <= to_signed(0,14);
 taps(274) <= to_signed(0,14);
 taps(275) <= to_signed(0,14);
 taps(276) <= to_signed(0,14);
 taps(277) <= to_signed(0,14);
 taps(278) <= to_signed(0,14);
 taps(279) <= to_signed(0,14);
 taps(280) <= to_signed(0,14);
 taps(281) <= to_signed(0,14);
 taps(282) <= to_signed(0,14);
 taps(283) <= to_signed(0,14);
 taps(284) <= to_signed(0,14);
 taps(285) <= to_signed(0,14);
 taps(286) <= to_signed(0,14);
 taps(287) <= to_signed(0,14);
 taps(288) <= to_signed(0,14);
 taps(289) <= to_signed(0,14);
 taps(290) <= to_signed(0,14);
 taps(291) <= to_signed(0,14);
 taps(292) <= to_signed(0,14);
 taps(293) <= to_signed(0,14);
 taps(294) <= to_signed(0,14);
 taps(295) <= to_signed(0,14);
 taps(296) <= to_signed(0,14);
 taps(297) <= to_signed(0,14);
 taps(298) <= to_signed(0,14);
 taps(299) <= to_signed(0,14);
 taps(300) <= to_signed(0,14);
 taps(301) <= to_signed(0,14);
 taps(302) <= to_signed(0,14);
 taps(303) <= to_signed(0,14);
 taps(304) <= to_signed(0,14);
 taps(305) <= to_signed(0,14);
 taps(306) <= to_signed(0,14);
 taps(307) <= to_signed(0,14);
 taps(308) <= to_signed(0,14);
 taps(309) <= to_signed(0,14);
 taps(310) <= to_signed(0,14);
 taps(311) <= to_signed(0,14);
 taps(312) <= to_signed(0,14);
 taps(313) <= to_signed(0,14);
 taps(314) <= to_signed(0,14);
 taps(315) <= to_signed(0,14);
 taps(316) <= to_signed(0,14);
 taps(317) <= to_signed(0,14);
 taps(318) <= to_signed(0,14);
 taps(319) <= to_signed(0,14);
 taps(320) <= to_signed(0,14);
 taps(321) <= to_signed(0,14);
 taps(322) <= to_signed(0,14);
 taps(323) <= to_signed(0,14);
 taps(324) <= to_signed(0,14);
 taps(325) <= to_signed(0,14);
 taps(326) <= to_signed(0,14);
 taps(327) <= to_signed(0,14);
 taps(328) <= to_signed(0,14);
 taps(329) <= to_signed(0,14);
 taps(330) <= to_signed(0,14);
 taps(331) <= to_signed(0,14);
 taps(332) <= to_signed(0,14);
 taps(333) <= to_signed(0,14);
 taps(334) <= to_signed(0,14);
 taps(335) <= to_signed(0,14);
 taps(336) <= to_signed(0,14);
 taps(337) <= to_signed(0,14);
 taps(338) <= to_signed(0,14);
 taps(339) <= to_signed(0,14);
 taps(340) <= to_signed(0,14);
 taps(341) <= to_signed(0,14);
 taps(342) <= to_signed(0,14);
 taps(343) <= to_signed(0,14);
 taps(344) <= to_signed(0,14);
 taps(345) <= to_signed(0,14);
 taps(346) <= to_signed(0,14);
 taps(347) <= to_signed(0,14);
 taps(348) <= to_signed(0,14);
 taps(349) <= to_signed(0,14);
 taps(350) <= to_signed(0,14);
 taps(351) <= to_signed(0,14);
 taps(352) <= to_signed(0,14);
 taps(353) <= to_signed(0,14);
 taps(354) <= to_signed(0,14);
 taps(355) <= to_signed(0,14);
 taps(356) <= to_signed(0,14);
 taps(357) <= to_signed(0,14);
 taps(358) <= to_signed(0,14);
 taps(359) <= to_signed(1,14);
 taps(360) <= to_signed(0,14);
 taps(361) <= to_signed(0,14);
 taps(362) <= to_signed(0,14);
 taps(363) <= to_signed(0,14);
 taps(364) <= to_signed(0,14);
 taps(365) <= to_signed(0,14);
 taps(366) <= to_signed(0,14);
 taps(367) <= to_signed(-1,14);
 taps(368) <= to_signed(-1,14);
 taps(369) <= to_signed(0,14);
 taps(370) <= to_signed(0,14);
 taps(371) <= to_signed(0,14);
 taps(372) <= to_signed(0,14);
 taps(373) <= to_signed(0,14);
 taps(374) <= to_signed(0,14);
 taps(375) <= to_signed(0,14);
 taps(376) <= to_signed(1,14);
 taps(377) <= to_signed(1,14);
 taps(378) <= to_signed(0,14);
 taps(379) <= to_signed(0,14);
 taps(380) <= to_signed(0,14);
 taps(381) <= to_signed(0,14);
 taps(382) <= to_signed(0,14);
 taps(383) <= to_signed(0,14);
 taps(384) <= to_signed(0,14);
 taps(385) <= to_signed(-1,14);
 taps(386) <= to_signed(0,14);
 taps(387) <= to_signed(0,14);
 taps(388) <= to_signed(0,14);
 taps(389) <= to_signed(0,14);
 taps(390) <= to_signed(0,14);
 taps(391) <= to_signed(0,14);
 taps(392) <= to_signed(0,14);
 taps(393) <= to_signed(0,14);
 taps(394) <= to_signed(0,14);
 taps(395) <= to_signed(0,14);
 taps(396) <= to_signed(0,14);
 taps(397) <= to_signed(0,14);
 taps(398) <= to_signed(0,14);
 taps(399) <= to_signed(0,14);
 taps(400) <= to_signed(0,14);
 taps(401) <= to_signed(0,14);
 taps(402) <= to_signed(0,14);
 taps(403) <= to_signed(0,14);
 taps(404) <= to_signed(0,14);
 taps(405) <= to_signed(0,14);
 taps(406) <= to_signed(0,14);
 taps(407) <= to_signed(0,14);
 taps(408) <= to_signed(0,14);
 taps(409) <= to_signed(0,14);
 taps(410) <= to_signed(0,14);
 taps(411) <= to_signed(0,14);
 taps(412) <= to_signed(0,14);
 taps(413) <= to_signed(0,14);
 taps(414) <= to_signed(0,14);
 taps(415) <= to_signed(0,14);
 taps(416) <= to_signed(0,14);
 taps(417) <= to_signed(0,14);
 taps(418) <= to_signed(0,14);
 taps(419) <= to_signed(0,14);
 taps(420) <= to_signed(0,14);
 taps(421) <= to_signed(0,14);
 taps(422) <= to_signed(0,14);
 taps(423) <= to_signed(0,14);
 taps(424) <= to_signed(0,14);
 taps(425) <= to_signed(0,14);
 taps(426) <= to_signed(0,14);
 taps(427) <= to_signed(0,14);
 taps(428) <= to_signed(0,14);
 taps(429) <= to_signed(0,14);
 taps(430) <= to_signed(0,14);
 taps(431) <= to_signed(0,14);
 taps(432) <= to_signed(0,14);
 taps(433) <= to_signed(0,14);
 taps(434) <= to_signed(0,14);
 taps(435) <= to_signed(0,14);
 taps(436) <= to_signed(0,14);
 taps(437) <= to_signed(1,14);
 taps(438) <= to_signed(1,14);
 taps(439) <= to_signed(0,14);
 taps(440) <= to_signed(0,14);
 taps(441) <= to_signed(0,14);
 taps(442) <= to_signed(0,14);
 taps(443) <= to_signed(0,14);
 taps(444) <= to_signed(-1,14);
 taps(445) <= to_signed(-1,14);
 taps(446) <= to_signed(-1,14);
 taps(447) <= to_signed(-1,14);
 taps(448) <= to_signed(-1,14);
 taps(449) <= to_signed(0,14);
 taps(450) <= to_signed(0,14);
 taps(451) <= to_signed(0,14);
 taps(452) <= to_signed(1,14);
 taps(453) <= to_signed(1,14);
 taps(454) <= to_signed(1,14);
 taps(455) <= to_signed(1,14);
 taps(456) <= to_signed(1,14);
 taps(457) <= to_signed(1,14);
 taps(458) <= to_signed(0,14);
 taps(459) <= to_signed(0,14);
 taps(460) <= to_signed(0,14);
 taps(461) <= to_signed(-1,14);
 taps(462) <= to_signed(-1,14);
 taps(463) <= to_signed(-1,14);
 taps(464) <= to_signed(-1,14);
 taps(465) <= to_signed(-1,14);
 taps(466) <= to_signed(-1,14);
 taps(467) <= to_signed(0,14);
 taps(468) <= to_signed(0,14);
 taps(469) <= to_signed(1,14);
 taps(470) <= to_signed(1,14);
 taps(471) <= to_signed(1,14);
 taps(472) <= to_signed(1,14);
 taps(473) <= to_signed(1,14);
 taps(474) <= to_signed(1,14);
 taps(475) <= to_signed(0,14);
 taps(476) <= to_signed(0,14);
 taps(477) <= to_signed(0,14);
 taps(478) <= to_signed(-1,14);
 taps(479) <= to_signed(-1,14);
 taps(480) <= to_signed(-1,14);
 taps(481) <= to_signed(-1,14);
 taps(482) <= to_signed(-1,14);
 taps(483) <= to_signed(-1,14);
 taps(484) <= to_signed(0,14);
 taps(485) <= to_signed(0,14);
 taps(486) <= to_signed(0,14);
 taps(487) <= to_signed(1,14);
 taps(488) <= to_signed(1,14);
 taps(489) <= to_signed(1,14);
 taps(490) <= to_signed(1,14);
 taps(491) <= to_signed(1,14);
 taps(492) <= to_signed(0,14);
 taps(493) <= to_signed(0,14);
 taps(494) <= to_signed(0,14);
 taps(495) <= to_signed(0,14);
 taps(496) <= to_signed(-1,14);
 taps(497) <= to_signed(-1,14);
 taps(498) <= to_signed(-1,14);
 taps(499) <= to_signed(-1,14);
 taps(500) <= to_signed(0,14);
 taps(501) <= to_signed(0,14);
 taps(502) <= to_signed(0,14);
 taps(503) <= to_signed(0,14);
 taps(504) <= to_signed(0,14);
 taps(505) <= to_signed(0,14);
 taps(506) <= to_signed(0,14);
 taps(507) <= to_signed(0,14);
 taps(508) <= to_signed(0,14);
 taps(509) <= to_signed(0,14);
 taps(510) <= to_signed(0,14);
 taps(511) <= to_signed(0,14);
 taps(512) <= to_signed(0,14);
 taps(513) <= to_signed(0,14);
 taps(514) <= to_signed(0,14);
 taps(515) <= to_signed(0,14);
 taps(516) <= to_signed(0,14);
 taps(517) <= to_signed(0,14);
 taps(518) <= to_signed(0,14);
 taps(519) <= to_signed(0,14);
 taps(520) <= to_signed(0,14);
 taps(521) <= to_signed(0,14);
 taps(522) <= to_signed(0,14);
 taps(523) <= to_signed(0,14);
 taps(524) <= to_signed(0,14);
 taps(525) <= to_signed(0,14);
 taps(526) <= to_signed(0,14);
 taps(527) <= to_signed(0,14);
 taps(528) <= to_signed(0,14);
 taps(529) <= to_signed(0,14);
 taps(530) <= to_signed(0,14);
 taps(531) <= to_signed(0,14);
 taps(532) <= to_signed(1,14);
 taps(533) <= to_signed(1,14);
 taps(534) <= to_signed(1,14);
 taps(535) <= to_signed(1,14);
 taps(536) <= to_signed(0,14);
 taps(537) <= to_signed(0,14);
 taps(538) <= to_signed(0,14);
 taps(539) <= to_signed(-1,14);
 taps(540) <= to_signed(-1,14);
 taps(541) <= to_signed(-1,14);
 taps(542) <= to_signed(-1,14);
 taps(543) <= to_signed(-1,14);
 taps(544) <= to_signed(-1,14);
 taps(545) <= to_signed(0,14);
 taps(546) <= to_signed(0,14);
 taps(547) <= to_signed(1,14);
 taps(548) <= to_signed(1,14);
 taps(549) <= to_signed(1,14);
 taps(550) <= to_signed(2,14);
 taps(551) <= to_signed(1,14);
 taps(552) <= to_signed(1,14);
 taps(553) <= to_signed(1,14);
 taps(554) <= to_signed(0,14);
 taps(555) <= to_signed(0,14);
 taps(556) <= to_signed(-1,14);
 taps(557) <= to_signed(-1,14);
 taps(558) <= to_signed(-2,14);
 taps(559) <= to_signed(-2,14);
 taps(560) <= to_signed(-2,14);
 taps(561) <= to_signed(-1,14);
 taps(562) <= to_signed(-1,14);
 taps(563) <= to_signed(0,14);
 taps(564) <= to_signed(1,14);
 taps(565) <= to_signed(1,14);
 taps(566) <= to_signed(2,14);
 taps(567) <= to_signed(2,14);
 taps(568) <= to_signed(2,14);
 taps(569) <= to_signed(2,14);
 taps(570) <= to_signed(1,14);
 taps(571) <= to_signed(1,14);
 taps(572) <= to_signed(0,14);
 taps(573) <= to_signed(-1,14);
 taps(574) <= to_signed(-2,14);
 taps(575) <= to_signed(-2,14);
 taps(576) <= to_signed(-2,14);
 taps(577) <= to_signed(-2,14);
 taps(578) <= to_signed(-2,14);
 taps(579) <= to_signed(-1,14);
 taps(580) <= to_signed(0,14);
 taps(581) <= to_signed(0,14);
 taps(582) <= to_signed(1,14);
 taps(583) <= to_signed(2,14);
 taps(584) <= to_signed(2,14);
 taps(585) <= to_signed(2,14);
 taps(586) <= to_signed(2,14);
 taps(587) <= to_signed(1,14);
 taps(588) <= to_signed(1,14);
 taps(589) <= to_signed(0,14);
 taps(590) <= to_signed(-1,14);
 taps(591) <= to_signed(-1,14);
 taps(592) <= to_signed(-2,14);
 taps(593) <= to_signed(-2,14);
 taps(594) <= to_signed(-2,14);
 taps(595) <= to_signed(-1,14);
 taps(596) <= to_signed(-1,14);
 taps(597) <= to_signed(0,14);
 taps(598) <= to_signed(0,14);
 taps(599) <= to_signed(1,14);
 taps(600) <= to_signed(1,14);
 taps(601) <= to_signed(1,14);
 taps(602) <= to_signed(1,14);
 taps(603) <= to_signed(1,14);
 taps(604) <= to_signed(1,14);
 taps(605) <= to_signed(1,14);
 taps(606) <= to_signed(0,14);
 taps(607) <= to_signed(0,14);
 taps(608) <= to_signed(-1,14);
 taps(609) <= to_signed(-1,14);
 taps(610) <= to_signed(-1,14);
 taps(611) <= to_signed(-1,14);
 taps(612) <= to_signed(-1,14);
 taps(613) <= to_signed(0,14);
 taps(614) <= to_signed(0,14);
 taps(615) <= to_signed(0,14);
 taps(616) <= to_signed(0,14);
 taps(617) <= to_signed(0,14);
 taps(618) <= to_signed(0,14);
 taps(619) <= to_signed(0,14);
 taps(620) <= to_signed(0,14);
 taps(621) <= to_signed(0,14);
 taps(622) <= to_signed(0,14);
 taps(623) <= to_signed(0,14);
 taps(624) <= to_signed(0,14);
 taps(625) <= to_signed(0,14);
 taps(626) <= to_signed(0,14);
 taps(627) <= to_signed(1,14);
 taps(628) <= to_signed(1,14);
 taps(629) <= to_signed(1,14);
 taps(630) <= to_signed(1,14);
 taps(631) <= to_signed(1,14);
 taps(632) <= to_signed(0,14);
 taps(633) <= to_signed(0,14);
 taps(634) <= to_signed(-1,14);
 taps(635) <= to_signed(-1,14);
 taps(636) <= to_signed(-2,14);
 taps(637) <= to_signed(-2,14);
 taps(638) <= to_signed(-2,14);
 taps(639) <= to_signed(-1,14);
 taps(640) <= to_signed(-1,14);
 taps(641) <= to_signed(0,14);
 taps(642) <= to_signed(1,14);
 taps(643) <= to_signed(1,14);
 taps(644) <= to_signed(2,14);
 taps(645) <= to_signed(2,14);
 taps(646) <= to_signed(3,14);
 taps(647) <= to_signed(2,14);
 taps(648) <= to_signed(2,14);
 taps(649) <= to_signed(1,14);
 taps(650) <= to_signed(0,14);
 taps(651) <= to_signed(-1,14);
 taps(652) <= to_signed(-2,14);
 taps(653) <= to_signed(-3,14);
 taps(654) <= to_signed(-3,14);
 taps(655) <= to_signed(-3,14);
 taps(656) <= to_signed(-3,14);
 taps(657) <= to_signed(-2,14);
 taps(658) <= to_signed(-1,14);
 taps(659) <= to_signed(0,14);
 taps(660) <= to_signed(2,14);
 taps(661) <= to_signed(3,14);
 taps(662) <= to_signed(4,14);
 taps(663) <= to_signed(4,14);
 taps(664) <= to_signed(4,14);
 taps(665) <= to_signed(3,14);
 taps(666) <= to_signed(2,14);
 taps(667) <= to_signed(0,14);
 taps(668) <= to_signed(-1,14);
 taps(669) <= to_signed(-2,14);
 taps(670) <= to_signed(-3,14);
 taps(671) <= to_signed(-4,14);
 taps(672) <= to_signed(-4,14);
 taps(673) <= to_signed(-4,14);
 taps(674) <= to_signed(-3,14);
 taps(675) <= to_signed(-1,14);
 taps(676) <= to_signed(0,14);
 taps(677) <= to_signed(1,14);
 taps(678) <= to_signed(3,14);
 taps(679) <= to_signed(4,14);
 taps(680) <= to_signed(4,14);
 taps(681) <= to_signed(4,14);
 taps(682) <= to_signed(3,14);
 taps(683) <= to_signed(2,14);
 taps(684) <= to_signed(1,14);
 taps(685) <= to_signed(0,14);
 taps(686) <= to_signed(-2,14);
 taps(687) <= to_signed(-3,14);
 taps(688) <= to_signed(-4,14);
 taps(689) <= to_signed(-4,14);
 taps(690) <= to_signed(-4,14);
 taps(691) <= to_signed(-3,14);
 taps(692) <= to_signed(-2,14);
 taps(693) <= to_signed(0,14);
 taps(694) <= to_signed(1,14);
 taps(695) <= to_signed(2,14);
 taps(696) <= to_signed(3,14);
 taps(697) <= to_signed(3,14);
 taps(698) <= to_signed(3,14);
 taps(699) <= to_signed(3,14);
 taps(700) <= to_signed(2,14);
 taps(701) <= to_signed(1,14);
 taps(702) <= to_signed(0,14);
 taps(703) <= to_signed(-1,14);
 taps(704) <= to_signed(-2,14);
 taps(705) <= to_signed(-2,14);
 taps(706) <= to_signed(-2,14);
 taps(707) <= to_signed(-2,14);
 taps(708) <= to_signed(-2,14);
 taps(709) <= to_signed(-1,14);
 taps(710) <= to_signed(0,14);
 taps(711) <= to_signed(0,14);
 taps(712) <= to_signed(1,14);
 taps(713) <= to_signed(1,14);
 taps(714) <= to_signed(1,14);
 taps(715) <= to_signed(1,14);
 taps(716) <= to_signed(1,14);
 taps(717) <= to_signed(0,14);
 taps(718) <= to_signed(0,14);
 taps(719) <= to_signed(0,14);
 taps(720) <= to_signed(0,14);
 taps(721) <= to_signed(0,14);
 taps(722) <= to_signed(0,14);
 taps(723) <= to_signed(1,14);
 taps(724) <= to_signed(1,14);
 taps(725) <= to_signed(1,14);
 taps(726) <= to_signed(1,14);
 taps(727) <= to_signed(1,14);
 taps(728) <= to_signed(0,14);
 taps(729) <= to_signed(0,14);
 taps(730) <= to_signed(-1,14);
 taps(731) <= to_signed(-2,14);
 taps(732) <= to_signed(-2,14);
 taps(733) <= to_signed(-3,14);
 taps(734) <= to_signed(-2,14);
 taps(735) <= to_signed(-2,14);
 taps(736) <= to_signed(-1,14);
 taps(737) <= to_signed(0,14);
 taps(738) <= to_signed(1,14);
 taps(739) <= to_signed(3,14);
 taps(740) <= to_signed(4,14);
 taps(741) <= to_signed(4,14);
 taps(742) <= to_signed(4,14);
 taps(743) <= to_signed(4,14);
 taps(744) <= to_signed(3,14);
 taps(745) <= to_signed(1,14);
 taps(746) <= to_signed(-1,14);
 taps(747) <= to_signed(-3,14);
 taps(748) <= to_signed(-4,14);
 taps(749) <= to_signed(-6,14);
 taps(750) <= to_signed(-6,14);
 taps(751) <= to_signed(-6,14);
 taps(752) <= to_signed(-5,14);
 taps(753) <= to_signed(-3,14);
 taps(754) <= to_signed(-1,14);
 taps(755) <= to_signed(2,14);
 taps(756) <= to_signed(4,14);
 taps(757) <= to_signed(6,14);
 taps(758) <= to_signed(7,14);
 taps(759) <= to_signed(8,14);
 taps(760) <= to_signed(7,14);
 taps(761) <= to_signed(5,14);
 taps(762) <= to_signed(3,14);
 taps(763) <= to_signed(0,14);
 taps(764) <= to_signed(-3,14);
 taps(765) <= to_signed(-6,14);
 taps(766) <= to_signed(-8,14);
 taps(767) <= to_signed(-9,14);
 taps(768) <= to_signed(-9,14);
 taps(769) <= to_signed(-7,14);
 taps(770) <= to_signed(-5,14);
 taps(771) <= to_signed(-2,14);
 taps(772) <= to_signed(1,14);
 taps(773) <= to_signed(5,14);
 taps(774) <= to_signed(7,14);
 taps(775) <= to_signed(9,14);
 taps(776) <= to_signed(9,14);
 taps(777) <= to_signed(9,14);
 taps(778) <= to_signed(7,14);
 taps(779) <= to_signed(4,14);
 taps(780) <= to_signed(1,14);
 taps(781) <= to_signed(-3,14);
 taps(782) <= to_signed(-6,14);
 taps(783) <= to_signed(-8,14);
 taps(784) <= to_signed(-9,14);
 taps(785) <= to_signed(-9,14);
 taps(786) <= to_signed(-8,14);
 taps(787) <= to_signed(-6,14);
 taps(788) <= to_signed(-3,14);
 taps(789) <= to_signed(0,14);
 taps(790) <= to_signed(3,14);
 taps(791) <= to_signed(6,14);
 taps(792) <= to_signed(8,14);
 taps(793) <= to_signed(9,14);
 taps(794) <= to_signed(8,14);
 taps(795) <= to_signed(7,14);
 taps(796) <= to_signed(5,14);
 taps(797) <= to_signed(2,14);
 taps(798) <= to_signed(-1,14);
 taps(799) <= to_signed(-4,14);
 taps(800) <= to_signed(-6,14);
 taps(801) <= to_signed(-7,14);
 taps(802) <= to_signed(-7,14);
 taps(803) <= to_signed(-6,14);
 taps(804) <= to_signed(-5,14);
 taps(805) <= to_signed(-3,14);
 taps(806) <= to_signed(-1,14);
 taps(807) <= to_signed(1,14);
 taps(808) <= to_signed(3,14);
 taps(809) <= to_signed(4,14);
 taps(810) <= to_signed(4,14);
 taps(811) <= to_signed(4,14);
 taps(812) <= to_signed(3,14);
 taps(813) <= to_signed(2,14);
 taps(814) <= to_signed(1,14);
 taps(815) <= to_signed(0,14);
 taps(816) <= to_signed(-1,14);
 taps(817) <= to_signed(-1,14);
 taps(818) <= to_signed(-1,14);
 taps(819) <= to_signed(-1,14);
 taps(820) <= to_signed(-1,14);
 taps(821) <= to_signed(0,14);
 taps(822) <= to_signed(0,14);
 taps(823) <= to_signed(0,14);
 taps(824) <= to_signed(0,14);
 taps(825) <= to_signed(-1,14);
 taps(826) <= to_signed(-2,14);
 taps(827) <= to_signed(-3,14);
 taps(828) <= to_signed(-3,14);
 taps(829) <= to_signed(-4,14);
 taps(830) <= to_signed(-3,14);
 taps(831) <= to_signed(-2,14);
 taps(832) <= to_signed(-1,14);
 taps(833) <= to_signed(1,14);
 taps(834) <= to_signed(4,14);
 taps(835) <= to_signed(6,14);
 taps(836) <= to_signed(8,14);
 taps(837) <= to_signed(8,14);
 taps(838) <= to_signed(8,14);
 taps(839) <= to_signed(7,14);
 taps(840) <= to_signed(4,14);
 taps(841) <= to_signed(0,14);
 taps(842) <= to_signed(-4,14);
 taps(843) <= to_signed(-8,14);
 taps(844) <= to_signed(-11,14);
 taps(845) <= to_signed(-13,14);
 taps(846) <= to_signed(-14,14);
 taps(847) <= to_signed(-12,14);
 taps(848) <= to_signed(-9,14);
 taps(849) <= to_signed(-4,14);
 taps(850) <= to_signed(1,14);
 taps(851) <= to_signed(7,14);
 taps(852) <= to_signed(13,14);
 taps(853) <= to_signed(17,14);
 taps(854) <= to_signed(19,14);
 taps(855) <= to_signed(18,14);
 taps(856) <= to_signed(15,14);
 taps(857) <= to_signed(10,14);
 taps(858) <= to_signed(3,14);
 taps(859) <= to_signed(-4,14);
 taps(860) <= to_signed(-12,14);
 taps(861) <= to_signed(-18,14);
 taps(862) <= to_signed(-22,14);
 taps(863) <= to_signed(-24,14);
 taps(864) <= to_signed(-22,14);
 taps(865) <= to_signed(-17,14);
 taps(866) <= to_signed(-10,14);
 taps(867) <= to_signed(-1,14);
 taps(868) <= to_signed(8,14);
 taps(869) <= to_signed(17,14);
 taps(870) <= to_signed(23,14);
 taps(871) <= to_signed(27,14);
 taps(872) <= to_signed(27,14);
 taps(873) <= to_signed(24,14);
 taps(874) <= to_signed(17,14);
 taps(875) <= to_signed(8,14);
 taps(876) <= to_signed(-2,14);
 taps(877) <= to_signed(-12,14);
 taps(878) <= to_signed(-21,14);
 taps(879) <= to_signed(-27,14);
 taps(880) <= to_signed(-30,14);
 taps(881) <= to_signed(-29,14);
 taps(882) <= to_signed(-24,14);
 taps(883) <= to_signed(-16,14);
 taps(884) <= to_signed(-6,14);
 taps(885) <= to_signed(6,14);
 taps(886) <= to_signed(16,14);
 taps(887) <= to_signed(24,14);
 taps(888) <= to_signed(29,14);
 taps(889) <= to_signed(31,14);
 taps(890) <= to_signed(28,14);
 taps(891) <= to_signed(22,14);
 taps(892) <= to_signed(13,14);
 taps(893) <= to_signed(2,14);
 taps(894) <= to_signed(-9,14);
 taps(895) <= to_signed(-18,14);
 taps(896) <= to_signed(-25,14);
 taps(897) <= to_signed(-28,14);
 taps(898) <= to_signed(-28,14);
 taps(899) <= to_signed(-24,14);
 taps(900) <= to_signed(-17,14);
 taps(901) <= to_signed(-8,14);
 taps(902) <= to_signed(1,14);
 taps(903) <= to_signed(10,14);
 taps(904) <= to_signed(17,14);
 taps(905) <= to_signed(22,14);
 taps(906) <= to_signed(23,14);
 taps(907) <= to_signed(21,14);
 taps(908) <= to_signed(17,14);
 taps(909) <= to_signed(11,14);
 taps(910) <= to_signed(4,14);
 taps(911) <= to_signed(-3,14);
 taps(912) <= to_signed(-8,14);
 taps(913) <= to_signed(-12,14);
 taps(914) <= to_signed(-13,14);
 taps(915) <= to_signed(-13,14);
 taps(916) <= to_signed(-10,14);
 taps(917) <= to_signed(-7,14);
 taps(918) <= to_signed(-3,14);
 taps(919) <= to_signed(0,14);
 taps(920) <= to_signed(1,14);
 taps(921) <= to_signed(2,14);
 taps(922) <= to_signed(1,14);
 taps(923) <= to_signed(-1,14);
 taps(924) <= to_signed(-3,14);
 taps(925) <= to_signed(-5,14);
 taps(926) <= to_signed(-5,14);
 taps(927) <= to_signed(-3,14);
 taps(928) <= to_signed(0,14);
 taps(929) <= to_signed(6,14);
 taps(930) <= to_signed(12,14);
 taps(931) <= to_signed(18,14);
 taps(932) <= to_signed(23,14);
 taps(933) <= to_signed(25,14);
 taps(934) <= to_signed(24,14);
 taps(935) <= to_signed(18,14);
 taps(936) <= to_signed(8,14);
 taps(937) <= to_signed(-5,14);
 taps(938) <= to_signed(-20,14);
 taps(939) <= to_signed(-35,14);
 taps(940) <= to_signed(-46,14);
 taps(941) <= to_signed(-53,14);
 taps(942) <= to_signed(-53,14);
 taps(943) <= to_signed(-45,14);
 taps(944) <= to_signed(-30,14);
 taps(945) <= to_signed(-8,14);
 taps(946) <= to_signed(18,14);
 taps(947) <= to_signed(45,14);
 taps(948) <= to_signed(69,14);
 taps(949) <= to_signed(86,14);
 taps(950) <= to_signed(92,14);
 taps(951) <= to_signed(87,14);
 taps(952) <= to_signed(69,14);
 taps(953) <= to_signed(39,14);
 taps(954) <= to_signed(0,14);
 taps(955) <= to_signed(-42,14);
 taps(956) <= to_signed(-83,14);
 taps(957) <= to_signed(-117,14);
 taps(958) <= to_signed(-138,14);
 taps(959) <= to_signed(-141,14);
 taps(960) <= to_signed(-126,14);
 taps(961) <= to_signed(-91,14);
 taps(962) <= to_signed(-41,14);
 taps(963) <= to_signed(19,14);
 taps(964) <= to_signed(83,14);
 taps(965) <= to_signed(140,14);
 taps(966) <= to_signed(183,14);
 taps(967) <= to_signed(205,14);
 taps(968) <= to_signed(201,14);
 taps(969) <= to_signed(169,14);
 taps(970) <= to_signed(111,14);
 taps(971) <= to_signed(33,14);
 taps(972) <= to_signed(-56,14);
 taps(973) <= to_signed(-145,14);
 taps(974) <= to_signed(-221,14);
 taps(975) <= to_signed(-274,14);
 taps(976) <= to_signed(-293,14);
 taps(977) <= to_signed(-274,14);
 taps(978) <= to_signed(-217,14);
 taps(979) <= to_signed(-124,14);
 taps(980) <= to_signed(-8,14);
 taps(981) <= to_signed(119,14);
 taps(982) <= to_signed(240,14);
 taps(983) <= to_signed(339,14);
 taps(984) <= to_signed(399,14);
 taps(985) <= to_signed(411,14);
 taps(986) <= to_signed(367,14);
 taps(987) <= to_signed(269,14);
 taps(988) <= to_signed(127,14);
 taps(989) <= to_signed(-44,14);
 taps(990) <= to_signed(-225,14);
 taps(991) <= to_signed(-390,14);
 taps(992) <= to_signed(-517,14);
 taps(993) <= to_signed(-584,14);
 taps(994) <= to_signed(-579,14);
 taps(995) <= to_signed(-493,14);
 taps(996) <= to_signed(-332,14);
 taps(997) <= to_signed(-110,14);
 taps(998) <= to_signed(148,14);
 taps(999) <= to_signed(412,14);
 taps(1000) <= to_signed(647,14);
 taps(1001) <= to_signed(818,14);
 taps(1002) <= to_signed(896,14);
 taps(1003) <= to_signed(858,14);
 taps(1004) <= to_signed(698,14);
 taps(1005) <= to_signed(422,14);
 taps(1006) <= to_signed(51,14);
 taps(1007) <= to_signed(-376,14);
 taps(1008) <= to_signed(-811,14);
 taps(1009) <= to_signed(-1198,14);
 taps(1010) <= to_signed(-1478,14);
 taps(1011) <= to_signed(-1596,14);
 taps(1012) <= to_signed(-1510,14);
 taps(1013) <= to_signed(-1189,14);
 taps(1014) <= to_signed(-627,14);
 taps(1015) <= to_signed(164,14);
 taps(1016) <= to_signed(1147,14);
 taps(1017) <= to_signed(2266,14);
 taps(1018) <= to_signed(3448,14);
 taps(1019) <= to_signed(4612,14);
 taps(1020) <= to_signed(5672,14);
 taps(1021) <= to_signed(6549,14);
 taps(1022) <= to_signed(7175,14);
 taps(1023) <= to_signed(7501,14);
 taps(1024) <= to_signed(7501,14);
 taps(1025) <= to_signed(7175,14);
 taps(1026) <= to_signed(6549,14);
 taps(1027) <= to_signed(5672,14);
 taps(1028) <= to_signed(4612,14);
 taps(1029) <= to_signed(3448,14);
 taps(1030) <= to_signed(2266,14);
 taps(1031) <= to_signed(1147,14);
 taps(1032) <= to_signed(164,14);
 taps(1033) <= to_signed(-627,14);
 taps(1034) <= to_signed(-1189,14);
 taps(1035) <= to_signed(-1510,14);
 taps(1036) <= to_signed(-1596,14);
 taps(1037) <= to_signed(-1478,14);
 taps(1038) <= to_signed(-1198,14);
 taps(1039) <= to_signed(-811,14);
 taps(1040) <= to_signed(-376,14);
 taps(1041) <= to_signed(51,14);
 taps(1042) <= to_signed(422,14);
 taps(1043) <= to_signed(698,14);
 taps(1044) <= to_signed(858,14);
 taps(1045) <= to_signed(896,14);
 taps(1046) <= to_signed(818,14);
 taps(1047) <= to_signed(647,14);
 taps(1048) <= to_signed(412,14);
 taps(1049) <= to_signed(148,14);
 taps(1050) <= to_signed(-110,14);
 taps(1051) <= to_signed(-332,14);
 taps(1052) <= to_signed(-493,14);
 taps(1053) <= to_signed(-579,14);
 taps(1054) <= to_signed(-584,14);
 taps(1055) <= to_signed(-517,14);
 taps(1056) <= to_signed(-390,14);
 taps(1057) <= to_signed(-225,14);
 taps(1058) <= to_signed(-44,14);
 taps(1059) <= to_signed(127,14);
 taps(1060) <= to_signed(269,14);
 taps(1061) <= to_signed(367,14);
 taps(1062) <= to_signed(411,14);
 taps(1063) <= to_signed(399,14);
 taps(1064) <= to_signed(339,14);
 taps(1065) <= to_signed(240,14);
 taps(1066) <= to_signed(119,14);
 taps(1067) <= to_signed(-8,14);
 taps(1068) <= to_signed(-124,14);
 taps(1069) <= to_signed(-217,14);
 taps(1070) <= to_signed(-274,14);
 taps(1071) <= to_signed(-293,14);
 taps(1072) <= to_signed(-274,14);
 taps(1073) <= to_signed(-221,14);
 taps(1074) <= to_signed(-145,14);
 taps(1075) <= to_signed(-56,14);
 taps(1076) <= to_signed(33,14);
 taps(1077) <= to_signed(111,14);
 taps(1078) <= to_signed(169,14);
 taps(1079) <= to_signed(201,14);
 taps(1080) <= to_signed(205,14);
 taps(1081) <= to_signed(183,14);
 taps(1082) <= to_signed(140,14);
 taps(1083) <= to_signed(83,14);
 taps(1084) <= to_signed(19,14);
 taps(1085) <= to_signed(-41,14);
 taps(1086) <= to_signed(-91,14);
 taps(1087) <= to_signed(-126,14);
 taps(1088) <= to_signed(-141,14);
 taps(1089) <= to_signed(-138,14);
 taps(1090) <= to_signed(-117,14);
 taps(1091) <= to_signed(-83,14);
 taps(1092) <= to_signed(-42,14);
 taps(1093) <= to_signed(0,14);
 taps(1094) <= to_signed(39,14);
 taps(1095) <= to_signed(69,14);
 taps(1096) <= to_signed(87,14);
 taps(1097) <= to_signed(92,14);
 taps(1098) <= to_signed(86,14);
 taps(1099) <= to_signed(69,14);
 taps(1100) <= to_signed(45,14);
 taps(1101) <= to_signed(18,14);
 taps(1102) <= to_signed(-8,14);
 taps(1103) <= to_signed(-30,14);
 taps(1104) <= to_signed(-45,14);
 taps(1105) <= to_signed(-53,14);
 taps(1106) <= to_signed(-53,14);
 taps(1107) <= to_signed(-46,14);
 taps(1108) <= to_signed(-35,14);
 taps(1109) <= to_signed(-20,14);
 taps(1110) <= to_signed(-5,14);
 taps(1111) <= to_signed(8,14);
 taps(1112) <= to_signed(18,14);
 taps(1113) <= to_signed(24,14);
 taps(1114) <= to_signed(25,14);
 taps(1115) <= to_signed(23,14);
 taps(1116) <= to_signed(18,14);
 taps(1117) <= to_signed(12,14);
 taps(1118) <= to_signed(6,14);
 taps(1119) <= to_signed(0,14);
 taps(1120) <= to_signed(-3,14);
 taps(1121) <= to_signed(-5,14);
 taps(1122) <= to_signed(-5,14);
 taps(1123) <= to_signed(-3,14);
 taps(1124) <= to_signed(-1,14);
 taps(1125) <= to_signed(1,14);
 taps(1126) <= to_signed(2,14);
 taps(1127) <= to_signed(1,14);
 taps(1128) <= to_signed(0,14);
 taps(1129) <= to_signed(-3,14);
 taps(1130) <= to_signed(-7,14);
 taps(1131) <= to_signed(-10,14);
 taps(1132) <= to_signed(-13,14);
 taps(1133) <= to_signed(-13,14);
 taps(1134) <= to_signed(-12,14);
 taps(1135) <= to_signed(-8,14);
 taps(1136) <= to_signed(-3,14);
 taps(1137) <= to_signed(4,14);
 taps(1138) <= to_signed(11,14);
 taps(1139) <= to_signed(17,14);
 taps(1140) <= to_signed(21,14);
 taps(1141) <= to_signed(23,14);
 taps(1142) <= to_signed(22,14);
 taps(1143) <= to_signed(17,14);
 taps(1144) <= to_signed(10,14);
 taps(1145) <= to_signed(1,14);
 taps(1146) <= to_signed(-8,14);
 taps(1147) <= to_signed(-17,14);
 taps(1148) <= to_signed(-24,14);
 taps(1149) <= to_signed(-28,14);
 taps(1150) <= to_signed(-28,14);
 taps(1151) <= to_signed(-25,14);
 taps(1152) <= to_signed(-18,14);
 taps(1153) <= to_signed(-9,14);
 taps(1154) <= to_signed(2,14);
 taps(1155) <= to_signed(13,14);
 taps(1156) <= to_signed(22,14);
 taps(1157) <= to_signed(28,14);
 taps(1158) <= to_signed(31,14);
 taps(1159) <= to_signed(29,14);
 taps(1160) <= to_signed(24,14);
 taps(1161) <= to_signed(16,14);
 taps(1162) <= to_signed(6,14);
 taps(1163) <= to_signed(-6,14);
 taps(1164) <= to_signed(-16,14);
 taps(1165) <= to_signed(-24,14);
 taps(1166) <= to_signed(-29,14);
 taps(1167) <= to_signed(-30,14);
 taps(1168) <= to_signed(-27,14);
 taps(1169) <= to_signed(-21,14);
 taps(1170) <= to_signed(-12,14);
 taps(1171) <= to_signed(-2,14);
 taps(1172) <= to_signed(8,14);
 taps(1173) <= to_signed(17,14);
 taps(1174) <= to_signed(24,14);
 taps(1175) <= to_signed(27,14);
 taps(1176) <= to_signed(27,14);
 taps(1177) <= to_signed(23,14);
 taps(1178) <= to_signed(17,14);
 taps(1179) <= to_signed(8,14);
 taps(1180) <= to_signed(-1,14);
 taps(1181) <= to_signed(-10,14);
 taps(1182) <= to_signed(-17,14);
 taps(1183) <= to_signed(-22,14);
 taps(1184) <= to_signed(-24,14);
 taps(1185) <= to_signed(-22,14);
 taps(1186) <= to_signed(-18,14);
 taps(1187) <= to_signed(-12,14);
 taps(1188) <= to_signed(-4,14);
 taps(1189) <= to_signed(3,14);
 taps(1190) <= to_signed(10,14);
 taps(1191) <= to_signed(15,14);
 taps(1192) <= to_signed(18,14);
 taps(1193) <= to_signed(19,14);
 taps(1194) <= to_signed(17,14);
 taps(1195) <= to_signed(13,14);
 taps(1196) <= to_signed(7,14);
 taps(1197) <= to_signed(1,14);
 taps(1198) <= to_signed(-4,14);
 taps(1199) <= to_signed(-9,14);
 taps(1200) <= to_signed(-12,14);
 taps(1201) <= to_signed(-14,14);
 taps(1202) <= to_signed(-13,14);
 taps(1203) <= to_signed(-11,14);
 taps(1204) <= to_signed(-8,14);
 taps(1205) <= to_signed(-4,14);
 taps(1206) <= to_signed(0,14);
 taps(1207) <= to_signed(4,14);
 taps(1208) <= to_signed(7,14);
 taps(1209) <= to_signed(8,14);
 taps(1210) <= to_signed(8,14);
 taps(1211) <= to_signed(8,14);
 taps(1212) <= to_signed(6,14);
 taps(1213) <= to_signed(4,14);
 taps(1214) <= to_signed(1,14);
 taps(1215) <= to_signed(-1,14);
 taps(1216) <= to_signed(-2,14);
 taps(1217) <= to_signed(-3,14);
 taps(1218) <= to_signed(-4,14);
 taps(1219) <= to_signed(-3,14);
 taps(1220) <= to_signed(-3,14);
 taps(1221) <= to_signed(-2,14);
 taps(1222) <= to_signed(-1,14);
 taps(1223) <= to_signed(0,14);
 taps(1224) <= to_signed(0,14);
 taps(1225) <= to_signed(0,14);
 taps(1226) <= to_signed(0,14);
 taps(1227) <= to_signed(-1,14);
 taps(1228) <= to_signed(-1,14);
 taps(1229) <= to_signed(-1,14);
 taps(1230) <= to_signed(-1,14);
 taps(1231) <= to_signed(-1,14);
 taps(1232) <= to_signed(0,14);
 taps(1233) <= to_signed(1,14);
 taps(1234) <= to_signed(2,14);
 taps(1235) <= to_signed(3,14);
 taps(1236) <= to_signed(4,14);
 taps(1237) <= to_signed(4,14);
 taps(1238) <= to_signed(4,14);
 taps(1239) <= to_signed(3,14);
 taps(1240) <= to_signed(1,14);
 taps(1241) <= to_signed(-1,14);
 taps(1242) <= to_signed(-3,14);
 taps(1243) <= to_signed(-5,14);
 taps(1244) <= to_signed(-6,14);
 taps(1245) <= to_signed(-7,14);
 taps(1246) <= to_signed(-7,14);
 taps(1247) <= to_signed(-6,14);
 taps(1248) <= to_signed(-4,14);
 taps(1249) <= to_signed(-1,14);
 taps(1250) <= to_signed(2,14);
 taps(1251) <= to_signed(5,14);
 taps(1252) <= to_signed(7,14);
 taps(1253) <= to_signed(8,14);
 taps(1254) <= to_signed(9,14);
 taps(1255) <= to_signed(8,14);
 taps(1256) <= to_signed(6,14);
 taps(1257) <= to_signed(3,14);
 taps(1258) <= to_signed(0,14);
 taps(1259) <= to_signed(-3,14);
 taps(1260) <= to_signed(-6,14);
 taps(1261) <= to_signed(-8,14);
 taps(1262) <= to_signed(-9,14);
 taps(1263) <= to_signed(-9,14);
 taps(1264) <= to_signed(-8,14);
 taps(1265) <= to_signed(-6,14);
 taps(1266) <= to_signed(-3,14);
 taps(1267) <= to_signed(1,14);
 taps(1268) <= to_signed(4,14);
 taps(1269) <= to_signed(7,14);
 taps(1270) <= to_signed(9,14);
 taps(1271) <= to_signed(9,14);
 taps(1272) <= to_signed(9,14);
 taps(1273) <= to_signed(7,14);
 taps(1274) <= to_signed(5,14);
 taps(1275) <= to_signed(1,14);
 taps(1276) <= to_signed(-2,14);
 taps(1277) <= to_signed(-5,14);
 taps(1278) <= to_signed(-7,14);
 taps(1279) <= to_signed(-9,14);
 taps(1280) <= to_signed(-9,14);
 taps(1281) <= to_signed(-8,14);
 taps(1282) <= to_signed(-6,14);
 taps(1283) <= to_signed(-3,14);
 taps(1284) <= to_signed(0,14);
 taps(1285) <= to_signed(3,14);
 taps(1286) <= to_signed(5,14);
 taps(1287) <= to_signed(7,14);
 taps(1288) <= to_signed(8,14);
 taps(1289) <= to_signed(7,14);
 taps(1290) <= to_signed(6,14);
 taps(1291) <= to_signed(4,14);
 taps(1292) <= to_signed(2,14);
 taps(1293) <= to_signed(-1,14);
 taps(1294) <= to_signed(-3,14);
 taps(1295) <= to_signed(-5,14);
 taps(1296) <= to_signed(-6,14);
 taps(1297) <= to_signed(-6,14);
 taps(1298) <= to_signed(-6,14);
 taps(1299) <= to_signed(-4,14);
 taps(1300) <= to_signed(-3,14);
 taps(1301) <= to_signed(-1,14);
 taps(1302) <= to_signed(1,14);
 taps(1303) <= to_signed(3,14);
 taps(1304) <= to_signed(4,14);
 taps(1305) <= to_signed(4,14);
 taps(1306) <= to_signed(4,14);
 taps(1307) <= to_signed(4,14);
 taps(1308) <= to_signed(3,14);
 taps(1309) <= to_signed(1,14);
 taps(1310) <= to_signed(0,14);
 taps(1311) <= to_signed(-1,14);
 taps(1312) <= to_signed(-2,14);
 taps(1313) <= to_signed(-2,14);
 taps(1314) <= to_signed(-3,14);
 taps(1315) <= to_signed(-2,14);
 taps(1316) <= to_signed(-2,14);
 taps(1317) <= to_signed(-1,14);
 taps(1318) <= to_signed(0,14);
 taps(1319) <= to_signed(0,14);
 taps(1320) <= to_signed(1,14);
 taps(1321) <= to_signed(1,14);
 taps(1322) <= to_signed(1,14);
 taps(1323) <= to_signed(1,14);
 taps(1324) <= to_signed(1,14);
 taps(1325) <= to_signed(0,14);
 taps(1326) <= to_signed(0,14);
 taps(1327) <= to_signed(0,14);
 taps(1328) <= to_signed(0,14);
 taps(1329) <= to_signed(0,14);
 taps(1330) <= to_signed(0,14);
 taps(1331) <= to_signed(1,14);
 taps(1332) <= to_signed(1,14);
 taps(1333) <= to_signed(1,14);
 taps(1334) <= to_signed(1,14);
 taps(1335) <= to_signed(1,14);
 taps(1336) <= to_signed(0,14);
 taps(1337) <= to_signed(0,14);
 taps(1338) <= to_signed(-1,14);
 taps(1339) <= to_signed(-2,14);
 taps(1340) <= to_signed(-2,14);
 taps(1341) <= to_signed(-2,14);
 taps(1342) <= to_signed(-2,14);
 taps(1343) <= to_signed(-2,14);
 taps(1344) <= to_signed(-1,14);
 taps(1345) <= to_signed(0,14);
 taps(1346) <= to_signed(1,14);
 taps(1347) <= to_signed(2,14);
 taps(1348) <= to_signed(3,14);
 taps(1349) <= to_signed(3,14);
 taps(1350) <= to_signed(3,14);
 taps(1351) <= to_signed(3,14);
 taps(1352) <= to_signed(2,14);
 taps(1353) <= to_signed(1,14);
 taps(1354) <= to_signed(0,14);
 taps(1355) <= to_signed(-2,14);
 taps(1356) <= to_signed(-3,14);
 taps(1357) <= to_signed(-4,14);
 taps(1358) <= to_signed(-4,14);
 taps(1359) <= to_signed(-4,14);
 taps(1360) <= to_signed(-3,14);
 taps(1361) <= to_signed(-2,14);
 taps(1362) <= to_signed(0,14);
 taps(1363) <= to_signed(1,14);
 taps(1364) <= to_signed(2,14);
 taps(1365) <= to_signed(3,14);
 taps(1366) <= to_signed(4,14);
 taps(1367) <= to_signed(4,14);
 taps(1368) <= to_signed(4,14);
 taps(1369) <= to_signed(3,14);
 taps(1370) <= to_signed(1,14);
 taps(1371) <= to_signed(0,14);
 taps(1372) <= to_signed(-1,14);
 taps(1373) <= to_signed(-3,14);
 taps(1374) <= to_signed(-4,14);
 taps(1375) <= to_signed(-4,14);
 taps(1376) <= to_signed(-4,14);
 taps(1377) <= to_signed(-3,14);
 taps(1378) <= to_signed(-2,14);
 taps(1379) <= to_signed(-1,14);
 taps(1380) <= to_signed(0,14);
 taps(1381) <= to_signed(2,14);
 taps(1382) <= to_signed(3,14);
 taps(1383) <= to_signed(4,14);
 taps(1384) <= to_signed(4,14);
 taps(1385) <= to_signed(4,14);
 taps(1386) <= to_signed(3,14);
 taps(1387) <= to_signed(2,14);
 taps(1388) <= to_signed(0,14);
 taps(1389) <= to_signed(-1,14);
 taps(1390) <= to_signed(-2,14);
 taps(1391) <= to_signed(-3,14);
 taps(1392) <= to_signed(-3,14);
 taps(1393) <= to_signed(-3,14);
 taps(1394) <= to_signed(-3,14);
 taps(1395) <= to_signed(-2,14);
 taps(1396) <= to_signed(-1,14);
 taps(1397) <= to_signed(0,14);
 taps(1398) <= to_signed(1,14);
 taps(1399) <= to_signed(2,14);
 taps(1400) <= to_signed(2,14);
 taps(1401) <= to_signed(3,14);
 taps(1402) <= to_signed(2,14);
 taps(1403) <= to_signed(2,14);
 taps(1404) <= to_signed(1,14);
 taps(1405) <= to_signed(1,14);
 taps(1406) <= to_signed(0,14);
 taps(1407) <= to_signed(-1,14);
 taps(1408) <= to_signed(-1,14);
 taps(1409) <= to_signed(-2,14);
 taps(1410) <= to_signed(-2,14);
 taps(1411) <= to_signed(-2,14);
 taps(1412) <= to_signed(-1,14);
 taps(1413) <= to_signed(-1,14);
 taps(1414) <= to_signed(0,14);
 taps(1415) <= to_signed(0,14);
 taps(1416) <= to_signed(1,14);
 taps(1417) <= to_signed(1,14);
 taps(1418) <= to_signed(1,14);
 taps(1419) <= to_signed(1,14);
 taps(1420) <= to_signed(1,14);
 taps(1421) <= to_signed(0,14);
 taps(1422) <= to_signed(0,14);
 taps(1423) <= to_signed(0,14);
 taps(1424) <= to_signed(0,14);
 taps(1425) <= to_signed(0,14);
 taps(1426) <= to_signed(0,14);
 taps(1427) <= to_signed(0,14);
 taps(1428) <= to_signed(0,14);
 taps(1429) <= to_signed(0,14);
 taps(1430) <= to_signed(0,14);
 taps(1431) <= to_signed(0,14);
 taps(1432) <= to_signed(0,14);
 taps(1433) <= to_signed(0,14);
 taps(1434) <= to_signed(0,14);
 taps(1435) <= to_signed(-1,14);
 taps(1436) <= to_signed(-1,14);
 taps(1437) <= to_signed(-1,14);
 taps(1438) <= to_signed(-1,14);
 taps(1439) <= to_signed(-1,14);
 taps(1440) <= to_signed(0,14);
 taps(1441) <= to_signed(0,14);
 taps(1442) <= to_signed(1,14);
 taps(1443) <= to_signed(1,14);
 taps(1444) <= to_signed(1,14);
 taps(1445) <= to_signed(1,14);
 taps(1446) <= to_signed(1,14);
 taps(1447) <= to_signed(1,14);
 taps(1448) <= to_signed(1,14);
 taps(1449) <= to_signed(0,14);
 taps(1450) <= to_signed(0,14);
 taps(1451) <= to_signed(-1,14);
 taps(1452) <= to_signed(-1,14);
 taps(1453) <= to_signed(-2,14);
 taps(1454) <= to_signed(-2,14);
 taps(1455) <= to_signed(-2,14);
 taps(1456) <= to_signed(-1,14);
 taps(1457) <= to_signed(-1,14);
 taps(1458) <= to_signed(0,14);
 taps(1459) <= to_signed(1,14);
 taps(1460) <= to_signed(1,14);
 taps(1461) <= to_signed(2,14);
 taps(1462) <= to_signed(2,14);
 taps(1463) <= to_signed(2,14);
 taps(1464) <= to_signed(2,14);
 taps(1465) <= to_signed(1,14);
 taps(1466) <= to_signed(0,14);
 taps(1467) <= to_signed(0,14);
 taps(1468) <= to_signed(-1,14);
 taps(1469) <= to_signed(-2,14);
 taps(1470) <= to_signed(-2,14);
 taps(1471) <= to_signed(-2,14);
 taps(1472) <= to_signed(-2,14);
 taps(1473) <= to_signed(-2,14);
 taps(1474) <= to_signed(-1,14);
 taps(1475) <= to_signed(0,14);
 taps(1476) <= to_signed(1,14);
 taps(1477) <= to_signed(1,14);
 taps(1478) <= to_signed(2,14);
 taps(1479) <= to_signed(2,14);
 taps(1480) <= to_signed(2,14);
 taps(1481) <= to_signed(2,14);
 taps(1482) <= to_signed(1,14);
 taps(1483) <= to_signed(1,14);
 taps(1484) <= to_signed(0,14);
 taps(1485) <= to_signed(-1,14);
 taps(1486) <= to_signed(-1,14);
 taps(1487) <= to_signed(-2,14);
 taps(1488) <= to_signed(-2,14);
 taps(1489) <= to_signed(-2,14);
 taps(1490) <= to_signed(-1,14);
 taps(1491) <= to_signed(-1,14);
 taps(1492) <= to_signed(0,14);
 taps(1493) <= to_signed(0,14);
 taps(1494) <= to_signed(1,14);
 taps(1495) <= to_signed(1,14);
 taps(1496) <= to_signed(1,14);
 taps(1497) <= to_signed(2,14);
 taps(1498) <= to_signed(1,14);
 taps(1499) <= to_signed(1,14);
 taps(1500) <= to_signed(1,14);
 taps(1501) <= to_signed(0,14);
 taps(1502) <= to_signed(0,14);
 taps(1503) <= to_signed(-1,14);
 taps(1504) <= to_signed(-1,14);
 taps(1505) <= to_signed(-1,14);
 taps(1506) <= to_signed(-1,14);
 taps(1507) <= to_signed(-1,14);
 taps(1508) <= to_signed(-1,14);
 taps(1509) <= to_signed(0,14);
 taps(1510) <= to_signed(0,14);
 taps(1511) <= to_signed(0,14);
 taps(1512) <= to_signed(1,14);
 taps(1513) <= to_signed(1,14);
 taps(1514) <= to_signed(1,14);
 taps(1515) <= to_signed(1,14);
 taps(1516) <= to_signed(0,14);
 taps(1517) <= to_signed(0,14);
 taps(1518) <= to_signed(0,14);
 taps(1519) <= to_signed(0,14);
 taps(1520) <= to_signed(0,14);
 taps(1521) <= to_signed(0,14);
 taps(1522) <= to_signed(0,14);
 taps(1523) <= to_signed(0,14);
 taps(1524) <= to_signed(0,14);
 taps(1525) <= to_signed(0,14);
 taps(1526) <= to_signed(0,14);
 taps(1527) <= to_signed(0,14);
 taps(1528) <= to_signed(0,14);
 taps(1529) <= to_signed(0,14);
 taps(1530) <= to_signed(0,14);
 taps(1531) <= to_signed(0,14);
 taps(1532) <= to_signed(0,14);
 taps(1533) <= to_signed(0,14);
 taps(1534) <= to_signed(0,14);
 taps(1535) <= to_signed(0,14);
 taps(1536) <= to_signed(0,14);
 taps(1537) <= to_signed(0,14);
 taps(1538) <= to_signed(0,14);
 taps(1539) <= to_signed(0,14);
 taps(1540) <= to_signed(0,14);
 taps(1541) <= to_signed(0,14);
 taps(1542) <= to_signed(0,14);
 taps(1543) <= to_signed(0,14);
 taps(1544) <= to_signed(0,14);
 taps(1545) <= to_signed(0,14);
 taps(1546) <= to_signed(0,14);
 taps(1547) <= to_signed(0,14);
 taps(1548) <= to_signed(-1,14);
 taps(1549) <= to_signed(-1,14);
 taps(1550) <= to_signed(-1,14);
 taps(1551) <= to_signed(-1,14);
 taps(1552) <= to_signed(0,14);
 taps(1553) <= to_signed(0,14);
 taps(1554) <= to_signed(0,14);
 taps(1555) <= to_signed(0,14);
 taps(1556) <= to_signed(1,14);
 taps(1557) <= to_signed(1,14);
 taps(1558) <= to_signed(1,14);
 taps(1559) <= to_signed(1,14);
 taps(1560) <= to_signed(1,14);
 taps(1561) <= to_signed(0,14);
 taps(1562) <= to_signed(0,14);
 taps(1563) <= to_signed(0,14);
 taps(1564) <= to_signed(-1,14);
 taps(1565) <= to_signed(-1,14);
 taps(1566) <= to_signed(-1,14);
 taps(1567) <= to_signed(-1,14);
 taps(1568) <= to_signed(-1,14);
 taps(1569) <= to_signed(-1,14);
 taps(1570) <= to_signed(0,14);
 taps(1571) <= to_signed(0,14);
 taps(1572) <= to_signed(0,14);
 taps(1573) <= to_signed(1,14);
 taps(1574) <= to_signed(1,14);
 taps(1575) <= to_signed(1,14);
 taps(1576) <= to_signed(1,14);
 taps(1577) <= to_signed(1,14);
 taps(1578) <= to_signed(1,14);
 taps(1579) <= to_signed(0,14);
 taps(1580) <= to_signed(0,14);
 taps(1581) <= to_signed(-1,14);
 taps(1582) <= to_signed(-1,14);
 taps(1583) <= to_signed(-1,14);
 taps(1584) <= to_signed(-1,14);
 taps(1585) <= to_signed(-1,14);
 taps(1586) <= to_signed(-1,14);
 taps(1587) <= to_signed(0,14);
 taps(1588) <= to_signed(0,14);
 taps(1589) <= to_signed(0,14);
 taps(1590) <= to_signed(1,14);
 taps(1591) <= to_signed(1,14);
 taps(1592) <= to_signed(1,14);
 taps(1593) <= to_signed(1,14);
 taps(1594) <= to_signed(1,14);
 taps(1595) <= to_signed(1,14);
 taps(1596) <= to_signed(0,14);
 taps(1597) <= to_signed(0,14);
 taps(1598) <= to_signed(0,14);
 taps(1599) <= to_signed(-1,14);
 taps(1600) <= to_signed(-1,14);
 taps(1601) <= to_signed(-1,14);
 taps(1602) <= to_signed(-1,14);
 taps(1603) <= to_signed(-1,14);
 taps(1604) <= to_signed(0,14);
 taps(1605) <= to_signed(0,14);
 taps(1606) <= to_signed(0,14);
 taps(1607) <= to_signed(0,14);
 taps(1608) <= to_signed(0,14);
 taps(1609) <= to_signed(1,14);
 taps(1610) <= to_signed(1,14);
 taps(1611) <= to_signed(0,14);
 taps(1612) <= to_signed(0,14);
 taps(1613) <= to_signed(0,14);
 taps(1614) <= to_signed(0,14);
 taps(1615) <= to_signed(0,14);
 taps(1616) <= to_signed(0,14);
 taps(1617) <= to_signed(0,14);
 taps(1618) <= to_signed(0,14);
 taps(1619) <= to_signed(0,14);
 taps(1620) <= to_signed(0,14);
 taps(1621) <= to_signed(0,14);
 taps(1622) <= to_signed(0,14);
 taps(1623) <= to_signed(0,14);
 taps(1624) <= to_signed(0,14);
 taps(1625) <= to_signed(0,14);
 taps(1626) <= to_signed(0,14);
 taps(1627) <= to_signed(0,14);
 taps(1628) <= to_signed(0,14);
 taps(1629) <= to_signed(0,14);
 taps(1630) <= to_signed(0,14);
 taps(1631) <= to_signed(0,14);
 taps(1632) <= to_signed(0,14);
 taps(1633) <= to_signed(0,14);
 taps(1634) <= to_signed(0,14);
 taps(1635) <= to_signed(0,14);
 taps(1636) <= to_signed(0,14);
 taps(1637) <= to_signed(0,14);
 taps(1638) <= to_signed(0,14);
 taps(1639) <= to_signed(0,14);
 taps(1640) <= to_signed(0,14);
 taps(1641) <= to_signed(0,14);
 taps(1642) <= to_signed(0,14);
 taps(1643) <= to_signed(0,14);
 taps(1644) <= to_signed(0,14);
 taps(1645) <= to_signed(0,14);
 taps(1646) <= to_signed(0,14);
 taps(1647) <= to_signed(0,14);
 taps(1648) <= to_signed(0,14);
 taps(1649) <= to_signed(0,14);
 taps(1650) <= to_signed(0,14);
 taps(1651) <= to_signed(0,14);
 taps(1652) <= to_signed(0,14);
 taps(1653) <= to_signed(0,14);
 taps(1654) <= to_signed(0,14);
 taps(1655) <= to_signed(0,14);
 taps(1656) <= to_signed(0,14);
 taps(1657) <= to_signed(0,14);
 taps(1658) <= to_signed(0,14);
 taps(1659) <= to_signed(0,14);
 taps(1660) <= to_signed(0,14);
 taps(1661) <= to_signed(0,14);
 taps(1662) <= to_signed(-1,14);
 taps(1663) <= to_signed(0,14);
 taps(1664) <= to_signed(0,14);
 taps(1665) <= to_signed(0,14);
 taps(1666) <= to_signed(0,14);
 taps(1667) <= to_signed(0,14);
 taps(1668) <= to_signed(0,14);
 taps(1669) <= to_signed(0,14);
 taps(1670) <= to_signed(1,14);
 taps(1671) <= to_signed(1,14);
 taps(1672) <= to_signed(0,14);
 taps(1673) <= to_signed(0,14);
 taps(1674) <= to_signed(0,14);
 taps(1675) <= to_signed(0,14);
 taps(1676) <= to_signed(0,14);
 taps(1677) <= to_signed(0,14);
 taps(1678) <= to_signed(0,14);
 taps(1679) <= to_signed(-1,14);
 taps(1680) <= to_signed(-1,14);
 taps(1681) <= to_signed(0,14);
 taps(1682) <= to_signed(0,14);
 taps(1683) <= to_signed(0,14);
 taps(1684) <= to_signed(0,14);
 taps(1685) <= to_signed(0,14);
 taps(1686) <= to_signed(0,14);
 taps(1687) <= to_signed(0,14);
 taps(1688) <= to_signed(1,14);
 taps(1689) <= to_signed(0,14);
 taps(1690) <= to_signed(0,14);
 taps(1691) <= to_signed(0,14);
 taps(1692) <= to_signed(0,14);
 taps(1693) <= to_signed(0,14);
 taps(1694) <= to_signed(0,14);
 taps(1695) <= to_signed(0,14);
 taps(1696) <= to_signed(0,14);
 taps(1697) <= to_signed(0,14);
 taps(1698) <= to_signed(0,14);
 taps(1699) <= to_signed(0,14);
 taps(1700) <= to_signed(0,14);
 taps(1701) <= to_signed(0,14);
 taps(1702) <= to_signed(0,14);
 taps(1703) <= to_signed(0,14);
 taps(1704) <= to_signed(0,14);
 taps(1705) <= to_signed(0,14);
 taps(1706) <= to_signed(0,14);
 taps(1707) <= to_signed(0,14);
 taps(1708) <= to_signed(0,14);
 taps(1709) <= to_signed(0,14);
 taps(1710) <= to_signed(0,14);
 taps(1711) <= to_signed(0,14);
 taps(1712) <= to_signed(0,14);
 taps(1713) <= to_signed(0,14);
 taps(1714) <= to_signed(0,14);
 taps(1715) <= to_signed(0,14);
 taps(1716) <= to_signed(0,14);
 taps(1717) <= to_signed(0,14);
 taps(1718) <= to_signed(0,14);
 taps(1719) <= to_signed(0,14);
 taps(1720) <= to_signed(0,14);
 taps(1721) <= to_signed(0,14);
 taps(1722) <= to_signed(0,14);
 taps(1723) <= to_signed(0,14);
 taps(1724) <= to_signed(0,14);
 taps(1725) <= to_signed(0,14);
 taps(1726) <= to_signed(0,14);
 taps(1727) <= to_signed(0,14);
 taps(1728) <= to_signed(0,14);
 taps(1729) <= to_signed(0,14);
 taps(1730) <= to_signed(0,14);
 taps(1731) <= to_signed(0,14);
 taps(1732) <= to_signed(0,14);
 taps(1733) <= to_signed(0,14);
 taps(1734) <= to_signed(0,14);
 taps(1735) <= to_signed(0,14);
 taps(1736) <= to_signed(0,14);
 taps(1737) <= to_signed(0,14);
 taps(1738) <= to_signed(0,14);
 taps(1739) <= to_signed(0,14);
 taps(1740) <= to_signed(0,14);
 taps(1741) <= to_signed(0,14);
 taps(1742) <= to_signed(0,14);
 taps(1743) <= to_signed(0,14);
 taps(1744) <= to_signed(0,14);
 taps(1745) <= to_signed(0,14);
 taps(1746) <= to_signed(0,14);
 taps(1747) <= to_signed(0,14);
 taps(1748) <= to_signed(0,14);
 taps(1749) <= to_signed(0,14);
 taps(1750) <= to_signed(0,14);
 taps(1751) <= to_signed(0,14);
 taps(1752) <= to_signed(0,14);
 taps(1753) <= to_signed(0,14);
 taps(1754) <= to_signed(0,14);
 taps(1755) <= to_signed(0,14);
 taps(1756) <= to_signed(0,14);
 taps(1757) <= to_signed(0,14);
 taps(1758) <= to_signed(0,14);
 taps(1759) <= to_signed(0,14);
 taps(1760) <= to_signed(0,14);
 taps(1761) <= to_signed(0,14);
 taps(1762) <= to_signed(0,14);
 taps(1763) <= to_signed(0,14);
 taps(1764) <= to_signed(0,14);
 taps(1765) <= to_signed(0,14);
 taps(1766) <= to_signed(0,14);
 taps(1767) <= to_signed(0,14);
 taps(1768) <= to_signed(0,14);
 taps(1769) <= to_signed(0,14);
 taps(1770) <= to_signed(0,14);
 taps(1771) <= to_signed(0,14);
 taps(1772) <= to_signed(0,14);
 taps(1773) <= to_signed(0,14);
 taps(1774) <= to_signed(0,14);
 taps(1775) <= to_signed(0,14);
 taps(1776) <= to_signed(0,14);
 taps(1777) <= to_signed(0,14);
 taps(1778) <= to_signed(0,14);
 taps(1779) <= to_signed(0,14);
 taps(1780) <= to_signed(0,14);
 taps(1781) <= to_signed(0,14);
 taps(1782) <= to_signed(0,14);
 taps(1783) <= to_signed(0,14);
 taps(1784) <= to_signed(0,14);
 taps(1785) <= to_signed(0,14);
 taps(1786) <= to_signed(0,14);
 taps(1787) <= to_signed(0,14);
 taps(1788) <= to_signed(0,14);
 taps(1789) <= to_signed(0,14);
 taps(1790) <= to_signed(0,14);
 taps(1791) <= to_signed(0,14);
 taps(1792) <= to_signed(0,14);
 taps(1793) <= to_signed(0,14);
 taps(1794) <= to_signed(0,14);
 taps(1795) <= to_signed(0,14);
 taps(1796) <= to_signed(0,14);
 taps(1797) <= to_signed(0,14);
 taps(1798) <= to_signed(0,14);
 taps(1799) <= to_signed(0,14);
 taps(1800) <= to_signed(0,14);
 taps(1801) <= to_signed(0,14);
 taps(1802) <= to_signed(0,14);
 taps(1803) <= to_signed(0,14);
 taps(1804) <= to_signed(0,14);
 taps(1805) <= to_signed(0,14);
 taps(1806) <= to_signed(0,14);
 taps(1807) <= to_signed(0,14);
 taps(1808) <= to_signed(0,14);
 taps(1809) <= to_signed(0,14);
 taps(1810) <= to_signed(0,14);
 taps(1811) <= to_signed(0,14);
 taps(1812) <= to_signed(0,14);
 taps(1813) <= to_signed(0,14);
 taps(1814) <= to_signed(0,14);
 taps(1815) <= to_signed(0,14);
 taps(1816) <= to_signed(0,14);
 taps(1817) <= to_signed(0,14);
 taps(1818) <= to_signed(0,14);
 taps(1819) <= to_signed(0,14);
 taps(1820) <= to_signed(0,14);
 taps(1821) <= to_signed(0,14);
 taps(1822) <= to_signed(0,14);
 taps(1823) <= to_signed(0,14);
 taps(1824) <= to_signed(0,14);
 taps(1825) <= to_signed(0,14);
 taps(1826) <= to_signed(0,14);
 taps(1827) <= to_signed(0,14);
 taps(1828) <= to_signed(0,14);
 taps(1829) <= to_signed(0,14);
 taps(1830) <= to_signed(0,14);
 taps(1831) <= to_signed(0,14);
 taps(1832) <= to_signed(0,14);
 taps(1833) <= to_signed(0,14);
 taps(1834) <= to_signed(0,14);
 taps(1835) <= to_signed(0,14);
 taps(1836) <= to_signed(0,14);
 taps(1837) <= to_signed(0,14);
 taps(1838) <= to_signed(0,14);
 taps(1839) <= to_signed(0,14);
 taps(1840) <= to_signed(0,14);
 taps(1841) <= to_signed(0,14);
 taps(1842) <= to_signed(0,14);
 taps(1843) <= to_signed(0,14);
 taps(1844) <= to_signed(0,14);
 taps(1845) <= to_signed(0,14);
 taps(1846) <= to_signed(0,14);
 taps(1847) <= to_signed(0,14);
 taps(1848) <= to_signed(0,14);
 taps(1849) <= to_signed(0,14);
 taps(1850) <= to_signed(0,14);
 taps(1851) <= to_signed(0,14);
 taps(1852) <= to_signed(0,14);
 taps(1853) <= to_signed(0,14);
 taps(1854) <= to_signed(0,14);
 taps(1855) <= to_signed(0,14);
 taps(1856) <= to_signed(0,14);
 taps(1857) <= to_signed(0,14);
 taps(1858) <= to_signed(0,14);
 taps(1859) <= to_signed(0,14);
 taps(1860) <= to_signed(0,14);
 taps(1861) <= to_signed(0,14);
 taps(1862) <= to_signed(0,14);
 taps(1863) <= to_signed(0,14);
 taps(1864) <= to_signed(0,14);
 taps(1865) <= to_signed(0,14);
 taps(1866) <= to_signed(0,14);
 taps(1867) <= to_signed(0,14);
 taps(1868) <= to_signed(0,14);
 taps(1869) <= to_signed(0,14);
 taps(1870) <= to_signed(0,14);
 taps(1871) <= to_signed(0,14);
 taps(1872) <= to_signed(0,14);
 taps(1873) <= to_signed(0,14);
 taps(1874) <= to_signed(0,14);
 taps(1875) <= to_signed(0,14);
 taps(1876) <= to_signed(0,14);
 taps(1877) <= to_signed(0,14);
 taps(1878) <= to_signed(0,14);
 taps(1879) <= to_signed(0,14);
 taps(1880) <= to_signed(0,14);
 taps(1881) <= to_signed(0,14);
 taps(1882) <= to_signed(0,14);
 taps(1883) <= to_signed(0,14);
 taps(1884) <= to_signed(0,14);
 taps(1885) <= to_signed(0,14);
 taps(1886) <= to_signed(0,14);
 taps(1887) <= to_signed(0,14);
 taps(1888) <= to_signed(0,14);
 taps(1889) <= to_signed(0,14);
 taps(1890) <= to_signed(0,14);
 taps(1891) <= to_signed(0,14);
 taps(1892) <= to_signed(0,14);
 taps(1893) <= to_signed(0,14);
 taps(1894) <= to_signed(0,14);
 taps(1895) <= to_signed(0,14);
 taps(1896) <= to_signed(0,14);
 taps(1897) <= to_signed(0,14);
 taps(1898) <= to_signed(0,14);
 taps(1899) <= to_signed(0,14);
 taps(1900) <= to_signed(0,14);
 taps(1901) <= to_signed(0,14);
 taps(1902) <= to_signed(0,14);
 taps(1903) <= to_signed(0,14);
 taps(1904) <= to_signed(0,14);
 taps(1905) <= to_signed(0,14);
 taps(1906) <= to_signed(0,14);
 taps(1907) <= to_signed(0,14);
 taps(1908) <= to_signed(0,14);
 taps(1909) <= to_signed(0,14);
 taps(1910) <= to_signed(0,14);
 taps(1911) <= to_signed(0,14);
 taps(1912) <= to_signed(0,14);
 taps(1913) <= to_signed(0,14);
 taps(1914) <= to_signed(0,14);
 taps(1915) <= to_signed(0,14);
 taps(1916) <= to_signed(0,14);
 taps(1917) <= to_signed(0,14);
 taps(1918) <= to_signed(0,14);
 taps(1919) <= to_signed(0,14);
 taps(1920) <= to_signed(0,14);
 taps(1921) <= to_signed(0,14);
 taps(1922) <= to_signed(0,14);
 taps(1923) <= to_signed(0,14);
 taps(1924) <= to_signed(0,14);
 taps(1925) <= to_signed(0,14);
 taps(1926) <= to_signed(0,14);
 taps(1927) <= to_signed(0,14);
 taps(1928) <= to_signed(0,14);
 taps(1929) <= to_signed(0,14);
 taps(1930) <= to_signed(0,14);
 taps(1931) <= to_signed(0,14);
 taps(1932) <= to_signed(0,14);
 taps(1933) <= to_signed(0,14);
 taps(1934) <= to_signed(0,14);
 taps(1935) <= to_signed(0,14);
 taps(1936) <= to_signed(0,14);
 taps(1937) <= to_signed(0,14);
 taps(1938) <= to_signed(0,14);
 taps(1939) <= to_signed(0,14);
 taps(1940) <= to_signed(0,14);
 taps(1941) <= to_signed(0,14);
 taps(1942) <= to_signed(0,14);
 taps(1943) <= to_signed(0,14);
 taps(1944) <= to_signed(0,14);
 taps(1945) <= to_signed(0,14);
 taps(1946) <= to_signed(0,14);
 taps(1947) <= to_signed(0,14);
 taps(1948) <= to_signed(0,14);
 taps(1949) <= to_signed(0,14);
 taps(1950) <= to_signed(0,14);
 taps(1951) <= to_signed(0,14);
 taps(1952) <= to_signed(0,14);
 taps(1953) <= to_signed(0,14);
 taps(1954) <= to_signed(0,14);
 taps(1955) <= to_signed(0,14);
 taps(1956) <= to_signed(0,14);
 taps(1957) <= to_signed(0,14);
 taps(1958) <= to_signed(0,14);
 taps(1959) <= to_signed(0,14);
 taps(1960) <= to_signed(0,14);
 taps(1961) <= to_signed(0,14);
 taps(1962) <= to_signed(0,14);
 taps(1963) <= to_signed(0,14);
 taps(1964) <= to_signed(0,14);
 taps(1965) <= to_signed(0,14);
 taps(1966) <= to_signed(0,14);
 taps(1967) <= to_signed(0,14);
 taps(1968) <= to_signed(0,14);
 taps(1969) <= to_signed(0,14);
 taps(1970) <= to_signed(0,14);
 taps(1971) <= to_signed(0,14);
 taps(1972) <= to_signed(0,14);
 taps(1973) <= to_signed(0,14);
 taps(1974) <= to_signed(0,14);
 taps(1975) <= to_signed(0,14);
 taps(1976) <= to_signed(0,14);
 taps(1977) <= to_signed(0,14);
 taps(1978) <= to_signed(0,14);
 taps(1979) <= to_signed(0,14);
 taps(1980) <= to_signed(0,14);
 taps(1981) <= to_signed(0,14);
 taps(1982) <= to_signed(0,14);
 taps(1983) <= to_signed(0,14);
 taps(1984) <= to_signed(0,14);
 taps(1985) <= to_signed(0,14);
 taps(1986) <= to_signed(0,14);
 taps(1987) <= to_signed(0,14);
 taps(1988) <= to_signed(0,14);
 taps(1989) <= to_signed(0,14);
 taps(1990) <= to_signed(0,14);
 taps(1991) <= to_signed(0,14);
 taps(1992) <= to_signed(0,14);
 taps(1993) <= to_signed(0,14);
 taps(1994) <= to_signed(0,14);
 taps(1995) <= to_signed(0,14);
 taps(1996) <= to_signed(0,14);
 taps(1997) <= to_signed(0,14);
 taps(1998) <= to_signed(0,14);
 taps(1999) <= to_signed(0,14);
 taps(2000) <= to_signed(0,14);
 taps(2001) <= to_signed(0,14);
 taps(2002) <= to_signed(0,14);
 taps(2003) <= to_signed(0,14);
 taps(2004) <= to_signed(0,14);
 taps(2005) <= to_signed(0,14);
 taps(2006) <= to_signed(0,14);
 taps(2007) <= to_signed(0,14);
 taps(2008) <= to_signed(0,14);
 taps(2009) <= to_signed(0,14);
 taps(2010) <= to_signed(0,14);
 taps(2011) <= to_signed(0,14);
 taps(2012) <= to_signed(0,14);
 taps(2013) <= to_signed(0,14);
 taps(2014) <= to_signed(0,14);
 taps(2015) <= to_signed(0,14);
 taps(2016) <= to_signed(0,14);
 taps(2017) <= to_signed(0,14);
 taps(2018) <= to_signed(0,14);
 taps(2019) <= to_signed(0,14);
 taps(2020) <= to_signed(0,14);
 taps(2021) <= to_signed(0,14);
 taps(2022) <= to_signed(0,14);
 taps(2023) <= to_signed(0,14);
 taps(2024) <= to_signed(0,14);
 taps(2025) <= to_signed(0,14);
 taps(2026) <= to_signed(0,14);
 taps(2027) <= to_signed(0,14);
 taps(2028) <= to_signed(0,14);
 taps(2029) <= to_signed(0,14);
 taps(2030) <= to_signed(0,14);
 taps(2031) <= to_signed(0,14);
 taps(2032) <= to_signed(0,14);
 taps(2033) <= to_signed(0,14);
 taps(2034) <= to_signed(0,14);
 taps(2035) <= to_signed(0,14);
 taps(2036) <= to_signed(0,14);
 taps(2037) <= to_signed(0,14);
 taps(2038) <= to_signed(0,14);
 taps(2039) <= to_signed(0,14);
 taps(2040) <= to_signed(0,14);
 taps(2041) <= to_signed(0,14);
 taps(2042) <= to_signed(0,14);
 taps(2043) <= to_signed(0,14);
 taps(2044) <= to_signed(0,14);
 taps(2045) <= to_signed(0,14);
 taps(2046) <= to_signed(0,14);
 taps(2047) <= to_signed(0,14);
                                                                                                         
                                                                                                         
                                                                                                         
 end rtl;                                                                                                
