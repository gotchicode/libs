library IEEE;                                                                 
use IEEE.std_logic_1164.all;                                                  
use IEEE.numeric_std.all;                                                     
                                                                              
entity sinus_rom is                                                                  
 port (                                                                       
            clk             : in std_logic;                                   
            addr_in         : in std_logic_vector(11 downto 0);               
            rd_en           : in std_logic;                                   
                                                                              
            data_out        : out std_logic_vector(15 downto 0);              
            data_out_en     : out std_logic                                   
 );                                                                           
end entity sinus_rom;                                                                
                                                                              
architecture rtl of sinus_rom is                                                     
                                                                              
type ROM_type is array (0 to 4095) of std_logic_vector(15 downto 0);            
signal ROM: ROM_type;                                                         
                                                                              
begin                                                                         
ROM(0) <= std_logic_vector(to_signed(0,16));
ROM(1) <= std_logic_vector(to_signed(2,16));
ROM(2) <= std_logic_vector(to_signed(3,16));
ROM(3) <= std_logic_vector(to_signed(5,16));
ROM(4) <= std_logic_vector(to_signed(6,16));
ROM(5) <= std_logic_vector(to_signed(8,16));
ROM(6) <= std_logic_vector(to_signed(9,16));
ROM(7) <= std_logic_vector(to_signed(11,16));
ROM(8) <= std_logic_vector(to_signed(13,16));
ROM(9) <= std_logic_vector(to_signed(14,16));
ROM(10) <= std_logic_vector(to_signed(16,16));
ROM(11) <= std_logic_vector(to_signed(17,16));
ROM(12) <= std_logic_vector(to_signed(19,16));
ROM(13) <= std_logic_vector(to_signed(20,16));
ROM(14) <= std_logic_vector(to_signed(22,16));
ROM(15) <= std_logic_vector(to_signed(24,16));
ROM(16) <= std_logic_vector(to_signed(25,16));
ROM(17) <= std_logic_vector(to_signed(27,16));
ROM(18) <= std_logic_vector(to_signed(28,16));
ROM(19) <= std_logic_vector(to_signed(30,16));
ROM(20) <= std_logic_vector(to_signed(31,16));
ROM(21) <= std_logic_vector(to_signed(33,16));
ROM(22) <= std_logic_vector(to_signed(35,16));
ROM(23) <= std_logic_vector(to_signed(36,16));
ROM(24) <= std_logic_vector(to_signed(38,16));
ROM(25) <= std_logic_vector(to_signed(39,16));
ROM(26) <= std_logic_vector(to_signed(41,16));
ROM(27) <= std_logic_vector(to_signed(42,16));
ROM(28) <= std_logic_vector(to_signed(44,16));
ROM(29) <= std_logic_vector(to_signed(46,16));
ROM(30) <= std_logic_vector(to_signed(47,16));
ROM(31) <= std_logic_vector(to_signed(49,16));
ROM(32) <= std_logic_vector(to_signed(50,16));
ROM(33) <= std_logic_vector(to_signed(52,16));
ROM(34) <= std_logic_vector(to_signed(53,16));
ROM(35) <= std_logic_vector(to_signed(55,16));
ROM(36) <= std_logic_vector(to_signed(57,16));
ROM(37) <= std_logic_vector(to_signed(58,16));
ROM(38) <= std_logic_vector(to_signed(60,16));
ROM(39) <= std_logic_vector(to_signed(61,16));
ROM(40) <= std_logic_vector(to_signed(63,16));
ROM(41) <= std_logic_vector(to_signed(64,16));
ROM(42) <= std_logic_vector(to_signed(66,16));
ROM(43) <= std_logic_vector(to_signed(67,16));
ROM(44) <= std_logic_vector(to_signed(69,16));
ROM(45) <= std_logic_vector(to_signed(71,16));
ROM(46) <= std_logic_vector(to_signed(72,16));
ROM(47) <= std_logic_vector(to_signed(74,16));
ROM(48) <= std_logic_vector(to_signed(75,16));
ROM(49) <= std_logic_vector(to_signed(77,16));
ROM(50) <= std_logic_vector(to_signed(78,16));
ROM(51) <= std_logic_vector(to_signed(80,16));
ROM(52) <= std_logic_vector(to_signed(82,16));
ROM(53) <= std_logic_vector(to_signed(83,16));
ROM(54) <= std_logic_vector(to_signed(85,16));
ROM(55) <= std_logic_vector(to_signed(86,16));
ROM(56) <= std_logic_vector(to_signed(88,16));
ROM(57) <= std_logic_vector(to_signed(89,16));
ROM(58) <= std_logic_vector(to_signed(91,16));
ROM(59) <= std_logic_vector(to_signed(93,16));
ROM(60) <= std_logic_vector(to_signed(94,16));
ROM(61) <= std_logic_vector(to_signed(96,16));
ROM(62) <= std_logic_vector(to_signed(97,16));
ROM(63) <= std_logic_vector(to_signed(99,16));
ROM(64) <= std_logic_vector(to_signed(100,16));
ROM(65) <= std_logic_vector(to_signed(102,16));
ROM(66) <= std_logic_vector(to_signed(103,16));
ROM(67) <= std_logic_vector(to_signed(105,16));
ROM(68) <= std_logic_vector(to_signed(107,16));
ROM(69) <= std_logic_vector(to_signed(108,16));
ROM(70) <= std_logic_vector(to_signed(110,16));
ROM(71) <= std_logic_vector(to_signed(111,16));
ROM(72) <= std_logic_vector(to_signed(113,16));
ROM(73) <= std_logic_vector(to_signed(114,16));
ROM(74) <= std_logic_vector(to_signed(116,16));
ROM(75) <= std_logic_vector(to_signed(118,16));
ROM(76) <= std_logic_vector(to_signed(119,16));
ROM(77) <= std_logic_vector(to_signed(121,16));
ROM(78) <= std_logic_vector(to_signed(122,16));
ROM(79) <= std_logic_vector(to_signed(124,16));
ROM(80) <= std_logic_vector(to_signed(125,16));
ROM(81) <= std_logic_vector(to_signed(127,16));
ROM(82) <= std_logic_vector(to_signed(128,16));
ROM(83) <= std_logic_vector(to_signed(130,16));
ROM(84) <= std_logic_vector(to_signed(132,16));
ROM(85) <= std_logic_vector(to_signed(133,16));
ROM(86) <= std_logic_vector(to_signed(135,16));
ROM(87) <= std_logic_vector(to_signed(136,16));
ROM(88) <= std_logic_vector(to_signed(138,16));
ROM(89) <= std_logic_vector(to_signed(139,16));
ROM(90) <= std_logic_vector(to_signed(141,16));
ROM(91) <= std_logic_vector(to_signed(142,16));
ROM(92) <= std_logic_vector(to_signed(144,16));
ROM(93) <= std_logic_vector(to_signed(146,16));
ROM(94) <= std_logic_vector(to_signed(147,16));
ROM(95) <= std_logic_vector(to_signed(149,16));
ROM(96) <= std_logic_vector(to_signed(150,16));
ROM(97) <= std_logic_vector(to_signed(152,16));
ROM(98) <= std_logic_vector(to_signed(153,16));
ROM(99) <= std_logic_vector(to_signed(155,16));
ROM(100) <= std_logic_vector(to_signed(156,16));
ROM(101) <= std_logic_vector(to_signed(158,16));
ROM(102) <= std_logic_vector(to_signed(160,16));
ROM(103) <= std_logic_vector(to_signed(161,16));
ROM(104) <= std_logic_vector(to_signed(163,16));
ROM(105) <= std_logic_vector(to_signed(164,16));
ROM(106) <= std_logic_vector(to_signed(166,16));
ROM(107) <= std_logic_vector(to_signed(167,16));
ROM(108) <= std_logic_vector(to_signed(169,16));
ROM(109) <= std_logic_vector(to_signed(170,16));
ROM(110) <= std_logic_vector(to_signed(172,16));
ROM(111) <= std_logic_vector(to_signed(174,16));
ROM(112) <= std_logic_vector(to_signed(175,16));
ROM(113) <= std_logic_vector(to_signed(177,16));
ROM(114) <= std_logic_vector(to_signed(178,16));
ROM(115) <= std_logic_vector(to_signed(180,16));
ROM(116) <= std_logic_vector(to_signed(181,16));
ROM(117) <= std_logic_vector(to_signed(183,16));
ROM(118) <= std_logic_vector(to_signed(184,16));
ROM(119) <= std_logic_vector(to_signed(186,16));
ROM(120) <= std_logic_vector(to_signed(187,16));
ROM(121) <= std_logic_vector(to_signed(189,16));
ROM(122) <= std_logic_vector(to_signed(191,16));
ROM(123) <= std_logic_vector(to_signed(192,16));
ROM(124) <= std_logic_vector(to_signed(194,16));
ROM(125) <= std_logic_vector(to_signed(195,16));
ROM(126) <= std_logic_vector(to_signed(197,16));
ROM(127) <= std_logic_vector(to_signed(198,16));
ROM(128) <= std_logic_vector(to_signed(200,16));
ROM(129) <= std_logic_vector(to_signed(201,16));
ROM(130) <= std_logic_vector(to_signed(203,16));
ROM(131) <= std_logic_vector(to_signed(204,16));
ROM(132) <= std_logic_vector(to_signed(206,16));
ROM(133) <= std_logic_vector(to_signed(207,16));
ROM(134) <= std_logic_vector(to_signed(209,16));
ROM(135) <= std_logic_vector(to_signed(211,16));
ROM(136) <= std_logic_vector(to_signed(212,16));
ROM(137) <= std_logic_vector(to_signed(214,16));
ROM(138) <= std_logic_vector(to_signed(215,16));
ROM(139) <= std_logic_vector(to_signed(217,16));
ROM(140) <= std_logic_vector(to_signed(218,16));
ROM(141) <= std_logic_vector(to_signed(220,16));
ROM(142) <= std_logic_vector(to_signed(221,16));
ROM(143) <= std_logic_vector(to_signed(223,16));
ROM(144) <= std_logic_vector(to_signed(224,16));
ROM(145) <= std_logic_vector(to_signed(226,16));
ROM(146) <= std_logic_vector(to_signed(227,16));
ROM(147) <= std_logic_vector(to_signed(229,16));
ROM(148) <= std_logic_vector(to_signed(230,16));
ROM(149) <= std_logic_vector(to_signed(232,16));
ROM(150) <= std_logic_vector(to_signed(234,16));
ROM(151) <= std_logic_vector(to_signed(235,16));
ROM(152) <= std_logic_vector(to_signed(237,16));
ROM(153) <= std_logic_vector(to_signed(238,16));
ROM(154) <= std_logic_vector(to_signed(240,16));
ROM(155) <= std_logic_vector(to_signed(241,16));
ROM(156) <= std_logic_vector(to_signed(243,16));
ROM(157) <= std_logic_vector(to_signed(244,16));
ROM(158) <= std_logic_vector(to_signed(246,16));
ROM(159) <= std_logic_vector(to_signed(247,16));
ROM(160) <= std_logic_vector(to_signed(249,16));
ROM(161) <= std_logic_vector(to_signed(250,16));
ROM(162) <= std_logic_vector(to_signed(252,16));
ROM(163) <= std_logic_vector(to_signed(253,16));
ROM(164) <= std_logic_vector(to_signed(255,16));
ROM(165) <= std_logic_vector(to_signed(256,16));
ROM(166) <= std_logic_vector(to_signed(258,16));
ROM(167) <= std_logic_vector(to_signed(259,16));
ROM(168) <= std_logic_vector(to_signed(261,16));
ROM(169) <= std_logic_vector(to_signed(263,16));
ROM(170) <= std_logic_vector(to_signed(264,16));
ROM(171) <= std_logic_vector(to_signed(266,16));
ROM(172) <= std_logic_vector(to_signed(267,16));
ROM(173) <= std_logic_vector(to_signed(269,16));
ROM(174) <= std_logic_vector(to_signed(270,16));
ROM(175) <= std_logic_vector(to_signed(272,16));
ROM(176) <= std_logic_vector(to_signed(273,16));
ROM(177) <= std_logic_vector(to_signed(275,16));
ROM(178) <= std_logic_vector(to_signed(276,16));
ROM(179) <= std_logic_vector(to_signed(278,16));
ROM(180) <= std_logic_vector(to_signed(279,16));
ROM(181) <= std_logic_vector(to_signed(281,16));
ROM(182) <= std_logic_vector(to_signed(282,16));
ROM(183) <= std_logic_vector(to_signed(284,16));
ROM(184) <= std_logic_vector(to_signed(285,16));
ROM(185) <= std_logic_vector(to_signed(287,16));
ROM(186) <= std_logic_vector(to_signed(288,16));
ROM(187) <= std_logic_vector(to_signed(290,16));
ROM(188) <= std_logic_vector(to_signed(291,16));
ROM(189) <= std_logic_vector(to_signed(293,16));
ROM(190) <= std_logic_vector(to_signed(294,16));
ROM(191) <= std_logic_vector(to_signed(296,16));
ROM(192) <= std_logic_vector(to_signed(297,16));
ROM(193) <= std_logic_vector(to_signed(299,16));
ROM(194) <= std_logic_vector(to_signed(300,16));
ROM(195) <= std_logic_vector(to_signed(302,16));
ROM(196) <= std_logic_vector(to_signed(303,16));
ROM(197) <= std_logic_vector(to_signed(305,16));
ROM(198) <= std_logic_vector(to_signed(306,16));
ROM(199) <= std_logic_vector(to_signed(308,16));
ROM(200) <= std_logic_vector(to_signed(309,16));
ROM(201) <= std_logic_vector(to_signed(311,16));
ROM(202) <= std_logic_vector(to_signed(312,16));
ROM(203) <= std_logic_vector(to_signed(314,16));
ROM(204) <= std_logic_vector(to_signed(315,16));
ROM(205) <= std_logic_vector(to_signed(317,16));
ROM(206) <= std_logic_vector(to_signed(318,16));
ROM(207) <= std_logic_vector(to_signed(320,16));
ROM(208) <= std_logic_vector(to_signed(321,16));
ROM(209) <= std_logic_vector(to_signed(323,16));
ROM(210) <= std_logic_vector(to_signed(324,16));
ROM(211) <= std_logic_vector(to_signed(326,16));
ROM(212) <= std_logic_vector(to_signed(327,16));
ROM(213) <= std_logic_vector(to_signed(329,16));
ROM(214) <= std_logic_vector(to_signed(330,16));
ROM(215) <= std_logic_vector(to_signed(332,16));
ROM(216) <= std_logic_vector(to_signed(333,16));
ROM(217) <= std_logic_vector(to_signed(335,16));
ROM(218) <= std_logic_vector(to_signed(336,16));
ROM(219) <= std_logic_vector(to_signed(338,16));
ROM(220) <= std_logic_vector(to_signed(339,16));
ROM(221) <= std_logic_vector(to_signed(341,16));
ROM(222) <= std_logic_vector(to_signed(342,16));
ROM(223) <= std_logic_vector(to_signed(343,16));
ROM(224) <= std_logic_vector(to_signed(345,16));
ROM(225) <= std_logic_vector(to_signed(346,16));
ROM(226) <= std_logic_vector(to_signed(348,16));
ROM(227) <= std_logic_vector(to_signed(349,16));
ROM(228) <= std_logic_vector(to_signed(351,16));
ROM(229) <= std_logic_vector(to_signed(352,16));
ROM(230) <= std_logic_vector(to_signed(354,16));
ROM(231) <= std_logic_vector(to_signed(355,16));
ROM(232) <= std_logic_vector(to_signed(357,16));
ROM(233) <= std_logic_vector(to_signed(358,16));
ROM(234) <= std_logic_vector(to_signed(360,16));
ROM(235) <= std_logic_vector(to_signed(361,16));
ROM(236) <= std_logic_vector(to_signed(363,16));
ROM(237) <= std_logic_vector(to_signed(364,16));
ROM(238) <= std_logic_vector(to_signed(366,16));
ROM(239) <= std_logic_vector(to_signed(367,16));
ROM(240) <= std_logic_vector(to_signed(369,16));
ROM(241) <= std_logic_vector(to_signed(370,16));
ROM(242) <= std_logic_vector(to_signed(371,16));
ROM(243) <= std_logic_vector(to_signed(373,16));
ROM(244) <= std_logic_vector(to_signed(374,16));
ROM(245) <= std_logic_vector(to_signed(376,16));
ROM(246) <= std_logic_vector(to_signed(377,16));
ROM(247) <= std_logic_vector(to_signed(379,16));
ROM(248) <= std_logic_vector(to_signed(380,16));
ROM(249) <= std_logic_vector(to_signed(382,16));
ROM(250) <= std_logic_vector(to_signed(383,16));
ROM(251) <= std_logic_vector(to_signed(385,16));
ROM(252) <= std_logic_vector(to_signed(386,16));
ROM(253) <= std_logic_vector(to_signed(388,16));
ROM(254) <= std_logic_vector(to_signed(389,16));
ROM(255) <= std_logic_vector(to_signed(390,16));
ROM(256) <= std_logic_vector(to_signed(392,16));
ROM(257) <= std_logic_vector(to_signed(393,16));
ROM(258) <= std_logic_vector(to_signed(395,16));
ROM(259) <= std_logic_vector(to_signed(396,16));
ROM(260) <= std_logic_vector(to_signed(398,16));
ROM(261) <= std_logic_vector(to_signed(399,16));
ROM(262) <= std_logic_vector(to_signed(401,16));
ROM(263) <= std_logic_vector(to_signed(402,16));
ROM(264) <= std_logic_vector(to_signed(403,16));
ROM(265) <= std_logic_vector(to_signed(405,16));
ROM(266) <= std_logic_vector(to_signed(406,16));
ROM(267) <= std_logic_vector(to_signed(408,16));
ROM(268) <= std_logic_vector(to_signed(409,16));
ROM(269) <= std_logic_vector(to_signed(411,16));
ROM(270) <= std_logic_vector(to_signed(412,16));
ROM(271) <= std_logic_vector(to_signed(414,16));
ROM(272) <= std_logic_vector(to_signed(415,16));
ROM(273) <= std_logic_vector(to_signed(416,16));
ROM(274) <= std_logic_vector(to_signed(418,16));
ROM(275) <= std_logic_vector(to_signed(419,16));
ROM(276) <= std_logic_vector(to_signed(421,16));
ROM(277) <= std_logic_vector(to_signed(422,16));
ROM(278) <= std_logic_vector(to_signed(424,16));
ROM(279) <= std_logic_vector(to_signed(425,16));
ROM(280) <= std_logic_vector(to_signed(426,16));
ROM(281) <= std_logic_vector(to_signed(428,16));
ROM(282) <= std_logic_vector(to_signed(429,16));
ROM(283) <= std_logic_vector(to_signed(431,16));
ROM(284) <= std_logic_vector(to_signed(432,16));
ROM(285) <= std_logic_vector(to_signed(434,16));
ROM(286) <= std_logic_vector(to_signed(435,16));
ROM(287) <= std_logic_vector(to_signed(436,16));
ROM(288) <= std_logic_vector(to_signed(438,16));
ROM(289) <= std_logic_vector(to_signed(439,16));
ROM(290) <= std_logic_vector(to_signed(441,16));
ROM(291) <= std_logic_vector(to_signed(442,16));
ROM(292) <= std_logic_vector(to_signed(443,16));
ROM(293) <= std_logic_vector(to_signed(445,16));
ROM(294) <= std_logic_vector(to_signed(446,16));
ROM(295) <= std_logic_vector(to_signed(448,16));
ROM(296) <= std_logic_vector(to_signed(449,16));
ROM(297) <= std_logic_vector(to_signed(451,16));
ROM(298) <= std_logic_vector(to_signed(452,16));
ROM(299) <= std_logic_vector(to_signed(453,16));
ROM(300) <= std_logic_vector(to_signed(455,16));
ROM(301) <= std_logic_vector(to_signed(456,16));
ROM(302) <= std_logic_vector(to_signed(458,16));
ROM(303) <= std_logic_vector(to_signed(459,16));
ROM(304) <= std_logic_vector(to_signed(460,16));
ROM(305) <= std_logic_vector(to_signed(462,16));
ROM(306) <= std_logic_vector(to_signed(463,16));
ROM(307) <= std_logic_vector(to_signed(465,16));
ROM(308) <= std_logic_vector(to_signed(466,16));
ROM(309) <= std_logic_vector(to_signed(467,16));
ROM(310) <= std_logic_vector(to_signed(469,16));
ROM(311) <= std_logic_vector(to_signed(470,16));
ROM(312) <= std_logic_vector(to_signed(472,16));
ROM(313) <= std_logic_vector(to_signed(473,16));
ROM(314) <= std_logic_vector(to_signed(474,16));
ROM(315) <= std_logic_vector(to_signed(476,16));
ROM(316) <= std_logic_vector(to_signed(477,16));
ROM(317) <= std_logic_vector(to_signed(479,16));
ROM(318) <= std_logic_vector(to_signed(480,16));
ROM(319) <= std_logic_vector(to_signed(481,16));
ROM(320) <= std_logic_vector(to_signed(483,16));
ROM(321) <= std_logic_vector(to_signed(484,16));
ROM(322) <= std_logic_vector(to_signed(485,16));
ROM(323) <= std_logic_vector(to_signed(487,16));
ROM(324) <= std_logic_vector(to_signed(488,16));
ROM(325) <= std_logic_vector(to_signed(490,16));
ROM(326) <= std_logic_vector(to_signed(491,16));
ROM(327) <= std_logic_vector(to_signed(492,16));
ROM(328) <= std_logic_vector(to_signed(494,16));
ROM(329) <= std_logic_vector(to_signed(495,16));
ROM(330) <= std_logic_vector(to_signed(497,16));
ROM(331) <= std_logic_vector(to_signed(498,16));
ROM(332) <= std_logic_vector(to_signed(499,16));
ROM(333) <= std_logic_vector(to_signed(501,16));
ROM(334) <= std_logic_vector(to_signed(502,16));
ROM(335) <= std_logic_vector(to_signed(503,16));
ROM(336) <= std_logic_vector(to_signed(505,16));
ROM(337) <= std_logic_vector(to_signed(506,16));
ROM(338) <= std_logic_vector(to_signed(507,16));
ROM(339) <= std_logic_vector(to_signed(509,16));
ROM(340) <= std_logic_vector(to_signed(510,16));
ROM(341) <= std_logic_vector(to_signed(512,16));
ROM(342) <= std_logic_vector(to_signed(513,16));
ROM(343) <= std_logic_vector(to_signed(514,16));
ROM(344) <= std_logic_vector(to_signed(516,16));
ROM(345) <= std_logic_vector(to_signed(517,16));
ROM(346) <= std_logic_vector(to_signed(518,16));
ROM(347) <= std_logic_vector(to_signed(520,16));
ROM(348) <= std_logic_vector(to_signed(521,16));
ROM(349) <= std_logic_vector(to_signed(522,16));
ROM(350) <= std_logic_vector(to_signed(524,16));
ROM(351) <= std_logic_vector(to_signed(525,16));
ROM(352) <= std_logic_vector(to_signed(526,16));
ROM(353) <= std_logic_vector(to_signed(528,16));
ROM(354) <= std_logic_vector(to_signed(529,16));
ROM(355) <= std_logic_vector(to_signed(530,16));
ROM(356) <= std_logic_vector(to_signed(532,16));
ROM(357) <= std_logic_vector(to_signed(533,16));
ROM(358) <= std_logic_vector(to_signed(535,16));
ROM(359) <= std_logic_vector(to_signed(536,16));
ROM(360) <= std_logic_vector(to_signed(537,16));
ROM(361) <= std_logic_vector(to_signed(539,16));
ROM(362) <= std_logic_vector(to_signed(540,16));
ROM(363) <= std_logic_vector(to_signed(541,16));
ROM(364) <= std_logic_vector(to_signed(543,16));
ROM(365) <= std_logic_vector(to_signed(544,16));
ROM(366) <= std_logic_vector(to_signed(545,16));
ROM(367) <= std_logic_vector(to_signed(547,16));
ROM(368) <= std_logic_vector(to_signed(548,16));
ROM(369) <= std_logic_vector(to_signed(549,16));
ROM(370) <= std_logic_vector(to_signed(550,16));
ROM(371) <= std_logic_vector(to_signed(552,16));
ROM(372) <= std_logic_vector(to_signed(553,16));
ROM(373) <= std_logic_vector(to_signed(554,16));
ROM(374) <= std_logic_vector(to_signed(556,16));
ROM(375) <= std_logic_vector(to_signed(557,16));
ROM(376) <= std_logic_vector(to_signed(558,16));
ROM(377) <= std_logic_vector(to_signed(560,16));
ROM(378) <= std_logic_vector(to_signed(561,16));
ROM(379) <= std_logic_vector(to_signed(562,16));
ROM(380) <= std_logic_vector(to_signed(564,16));
ROM(381) <= std_logic_vector(to_signed(565,16));
ROM(382) <= std_logic_vector(to_signed(566,16));
ROM(383) <= std_logic_vector(to_signed(568,16));
ROM(384) <= std_logic_vector(to_signed(569,16));
ROM(385) <= std_logic_vector(to_signed(570,16));
ROM(386) <= std_logic_vector(to_signed(572,16));
ROM(387) <= std_logic_vector(to_signed(573,16));
ROM(388) <= std_logic_vector(to_signed(574,16));
ROM(389) <= std_logic_vector(to_signed(575,16));
ROM(390) <= std_logic_vector(to_signed(577,16));
ROM(391) <= std_logic_vector(to_signed(578,16));
ROM(392) <= std_logic_vector(to_signed(579,16));
ROM(393) <= std_logic_vector(to_signed(581,16));
ROM(394) <= std_logic_vector(to_signed(582,16));
ROM(395) <= std_logic_vector(to_signed(583,16));
ROM(396) <= std_logic_vector(to_signed(584,16));
ROM(397) <= std_logic_vector(to_signed(586,16));
ROM(398) <= std_logic_vector(to_signed(587,16));
ROM(399) <= std_logic_vector(to_signed(588,16));
ROM(400) <= std_logic_vector(to_signed(590,16));
ROM(401) <= std_logic_vector(to_signed(591,16));
ROM(402) <= std_logic_vector(to_signed(592,16));
ROM(403) <= std_logic_vector(to_signed(593,16));
ROM(404) <= std_logic_vector(to_signed(595,16));
ROM(405) <= std_logic_vector(to_signed(596,16));
ROM(406) <= std_logic_vector(to_signed(597,16));
ROM(407) <= std_logic_vector(to_signed(599,16));
ROM(408) <= std_logic_vector(to_signed(600,16));
ROM(409) <= std_logic_vector(to_signed(601,16));
ROM(410) <= std_logic_vector(to_signed(602,16));
ROM(411) <= std_logic_vector(to_signed(604,16));
ROM(412) <= std_logic_vector(to_signed(605,16));
ROM(413) <= std_logic_vector(to_signed(606,16));
ROM(414) <= std_logic_vector(to_signed(607,16));
ROM(415) <= std_logic_vector(to_signed(609,16));
ROM(416) <= std_logic_vector(to_signed(610,16));
ROM(417) <= std_logic_vector(to_signed(611,16));
ROM(418) <= std_logic_vector(to_signed(613,16));
ROM(419) <= std_logic_vector(to_signed(614,16));
ROM(420) <= std_logic_vector(to_signed(615,16));
ROM(421) <= std_logic_vector(to_signed(616,16));
ROM(422) <= std_logic_vector(to_signed(618,16));
ROM(423) <= std_logic_vector(to_signed(619,16));
ROM(424) <= std_logic_vector(to_signed(620,16));
ROM(425) <= std_logic_vector(to_signed(621,16));
ROM(426) <= std_logic_vector(to_signed(623,16));
ROM(427) <= std_logic_vector(to_signed(624,16));
ROM(428) <= std_logic_vector(to_signed(625,16));
ROM(429) <= std_logic_vector(to_signed(626,16));
ROM(430) <= std_logic_vector(to_signed(628,16));
ROM(431) <= std_logic_vector(to_signed(629,16));
ROM(432) <= std_logic_vector(to_signed(630,16));
ROM(433) <= std_logic_vector(to_signed(631,16));
ROM(434) <= std_logic_vector(to_signed(632,16));
ROM(435) <= std_logic_vector(to_signed(634,16));
ROM(436) <= std_logic_vector(to_signed(635,16));
ROM(437) <= std_logic_vector(to_signed(636,16));
ROM(438) <= std_logic_vector(to_signed(637,16));
ROM(439) <= std_logic_vector(to_signed(639,16));
ROM(440) <= std_logic_vector(to_signed(640,16));
ROM(441) <= std_logic_vector(to_signed(641,16));
ROM(442) <= std_logic_vector(to_signed(642,16));
ROM(443) <= std_logic_vector(to_signed(644,16));
ROM(444) <= std_logic_vector(to_signed(645,16));
ROM(445) <= std_logic_vector(to_signed(646,16));
ROM(446) <= std_logic_vector(to_signed(647,16));
ROM(447) <= std_logic_vector(to_signed(648,16));
ROM(448) <= std_logic_vector(to_signed(650,16));
ROM(449) <= std_logic_vector(to_signed(651,16));
ROM(450) <= std_logic_vector(to_signed(652,16));
ROM(451) <= std_logic_vector(to_signed(653,16));
ROM(452) <= std_logic_vector(to_signed(654,16));
ROM(453) <= std_logic_vector(to_signed(656,16));
ROM(454) <= std_logic_vector(to_signed(657,16));
ROM(455) <= std_logic_vector(to_signed(658,16));
ROM(456) <= std_logic_vector(to_signed(659,16));
ROM(457) <= std_logic_vector(to_signed(660,16));
ROM(458) <= std_logic_vector(to_signed(662,16));
ROM(459) <= std_logic_vector(to_signed(663,16));
ROM(460) <= std_logic_vector(to_signed(664,16));
ROM(461) <= std_logic_vector(to_signed(665,16));
ROM(462) <= std_logic_vector(to_signed(666,16));
ROM(463) <= std_logic_vector(to_signed(668,16));
ROM(464) <= std_logic_vector(to_signed(669,16));
ROM(465) <= std_logic_vector(to_signed(670,16));
ROM(466) <= std_logic_vector(to_signed(671,16));
ROM(467) <= std_logic_vector(to_signed(672,16));
ROM(468) <= std_logic_vector(to_signed(674,16));
ROM(469) <= std_logic_vector(to_signed(675,16));
ROM(470) <= std_logic_vector(to_signed(676,16));
ROM(471) <= std_logic_vector(to_signed(677,16));
ROM(472) <= std_logic_vector(to_signed(678,16));
ROM(473) <= std_logic_vector(to_signed(679,16));
ROM(474) <= std_logic_vector(to_signed(681,16));
ROM(475) <= std_logic_vector(to_signed(682,16));
ROM(476) <= std_logic_vector(to_signed(683,16));
ROM(477) <= std_logic_vector(to_signed(684,16));
ROM(478) <= std_logic_vector(to_signed(685,16));
ROM(479) <= std_logic_vector(to_signed(687,16));
ROM(480) <= std_logic_vector(to_signed(688,16));
ROM(481) <= std_logic_vector(to_signed(689,16));
ROM(482) <= std_logic_vector(to_signed(690,16));
ROM(483) <= std_logic_vector(to_signed(691,16));
ROM(484) <= std_logic_vector(to_signed(692,16));
ROM(485) <= std_logic_vector(to_signed(693,16));
ROM(486) <= std_logic_vector(to_signed(695,16));
ROM(487) <= std_logic_vector(to_signed(696,16));
ROM(488) <= std_logic_vector(to_signed(697,16));
ROM(489) <= std_logic_vector(to_signed(698,16));
ROM(490) <= std_logic_vector(to_signed(699,16));
ROM(491) <= std_logic_vector(to_signed(700,16));
ROM(492) <= std_logic_vector(to_signed(702,16));
ROM(493) <= std_logic_vector(to_signed(703,16));
ROM(494) <= std_logic_vector(to_signed(704,16));
ROM(495) <= std_logic_vector(to_signed(705,16));
ROM(496) <= std_logic_vector(to_signed(706,16));
ROM(497) <= std_logic_vector(to_signed(707,16));
ROM(498) <= std_logic_vector(to_signed(708,16));
ROM(499) <= std_logic_vector(to_signed(709,16));
ROM(500) <= std_logic_vector(to_signed(711,16));
ROM(501) <= std_logic_vector(to_signed(712,16));
ROM(502) <= std_logic_vector(to_signed(713,16));
ROM(503) <= std_logic_vector(to_signed(714,16));
ROM(504) <= std_logic_vector(to_signed(715,16));
ROM(505) <= std_logic_vector(to_signed(716,16));
ROM(506) <= std_logic_vector(to_signed(717,16));
ROM(507) <= std_logic_vector(to_signed(719,16));
ROM(508) <= std_logic_vector(to_signed(720,16));
ROM(509) <= std_logic_vector(to_signed(721,16));
ROM(510) <= std_logic_vector(to_signed(722,16));
ROM(511) <= std_logic_vector(to_signed(723,16));
ROM(512) <= std_logic_vector(to_signed(724,16));
ROM(513) <= std_logic_vector(to_signed(725,16));
ROM(514) <= std_logic_vector(to_signed(726,16));
ROM(515) <= std_logic_vector(to_signed(727,16));
ROM(516) <= std_logic_vector(to_signed(729,16));
ROM(517) <= std_logic_vector(to_signed(730,16));
ROM(518) <= std_logic_vector(to_signed(731,16));
ROM(519) <= std_logic_vector(to_signed(732,16));
ROM(520) <= std_logic_vector(to_signed(733,16));
ROM(521) <= std_logic_vector(to_signed(734,16));
ROM(522) <= std_logic_vector(to_signed(735,16));
ROM(523) <= std_logic_vector(to_signed(736,16));
ROM(524) <= std_logic_vector(to_signed(737,16));
ROM(525) <= std_logic_vector(to_signed(738,16));
ROM(526) <= std_logic_vector(to_signed(739,16));
ROM(527) <= std_logic_vector(to_signed(741,16));
ROM(528) <= std_logic_vector(to_signed(742,16));
ROM(529) <= std_logic_vector(to_signed(743,16));
ROM(530) <= std_logic_vector(to_signed(744,16));
ROM(531) <= std_logic_vector(to_signed(745,16));
ROM(532) <= std_logic_vector(to_signed(746,16));
ROM(533) <= std_logic_vector(to_signed(747,16));
ROM(534) <= std_logic_vector(to_signed(748,16));
ROM(535) <= std_logic_vector(to_signed(749,16));
ROM(536) <= std_logic_vector(to_signed(750,16));
ROM(537) <= std_logic_vector(to_signed(751,16));
ROM(538) <= std_logic_vector(to_signed(752,16));
ROM(539) <= std_logic_vector(to_signed(753,16));
ROM(540) <= std_logic_vector(to_signed(755,16));
ROM(541) <= std_logic_vector(to_signed(756,16));
ROM(542) <= std_logic_vector(to_signed(757,16));
ROM(543) <= std_logic_vector(to_signed(758,16));
ROM(544) <= std_logic_vector(to_signed(759,16));
ROM(545) <= std_logic_vector(to_signed(760,16));
ROM(546) <= std_logic_vector(to_signed(761,16));
ROM(547) <= std_logic_vector(to_signed(762,16));
ROM(548) <= std_logic_vector(to_signed(763,16));
ROM(549) <= std_logic_vector(to_signed(764,16));
ROM(550) <= std_logic_vector(to_signed(765,16));
ROM(551) <= std_logic_vector(to_signed(766,16));
ROM(552) <= std_logic_vector(to_signed(767,16));
ROM(553) <= std_logic_vector(to_signed(768,16));
ROM(554) <= std_logic_vector(to_signed(769,16));
ROM(555) <= std_logic_vector(to_signed(770,16));
ROM(556) <= std_logic_vector(to_signed(771,16));
ROM(557) <= std_logic_vector(to_signed(772,16));
ROM(558) <= std_logic_vector(to_signed(773,16));
ROM(559) <= std_logic_vector(to_signed(774,16));
ROM(560) <= std_logic_vector(to_signed(775,16));
ROM(561) <= std_logic_vector(to_signed(776,16));
ROM(562) <= std_logic_vector(to_signed(777,16));
ROM(563) <= std_logic_vector(to_signed(778,16));
ROM(564) <= std_logic_vector(to_signed(779,16));
ROM(565) <= std_logic_vector(to_signed(780,16));
ROM(566) <= std_logic_vector(to_signed(782,16));
ROM(567) <= std_logic_vector(to_signed(783,16));
ROM(568) <= std_logic_vector(to_signed(784,16));
ROM(569) <= std_logic_vector(to_signed(785,16));
ROM(570) <= std_logic_vector(to_signed(786,16));
ROM(571) <= std_logic_vector(to_signed(787,16));
ROM(572) <= std_logic_vector(to_signed(788,16));
ROM(573) <= std_logic_vector(to_signed(789,16));
ROM(574) <= std_logic_vector(to_signed(790,16));
ROM(575) <= std_logic_vector(to_signed(791,16));
ROM(576) <= std_logic_vector(to_signed(792,16));
ROM(577) <= std_logic_vector(to_signed(793,16));
ROM(578) <= std_logic_vector(to_signed(794,16));
ROM(579) <= std_logic_vector(to_signed(795,16));
ROM(580) <= std_logic_vector(to_signed(796,16));
ROM(581) <= std_logic_vector(to_signed(797,16));
ROM(582) <= std_logic_vector(to_signed(798,16));
ROM(583) <= std_logic_vector(to_signed(798,16));
ROM(584) <= std_logic_vector(to_signed(799,16));
ROM(585) <= std_logic_vector(to_signed(800,16));
ROM(586) <= std_logic_vector(to_signed(801,16));
ROM(587) <= std_logic_vector(to_signed(802,16));
ROM(588) <= std_logic_vector(to_signed(803,16));
ROM(589) <= std_logic_vector(to_signed(804,16));
ROM(590) <= std_logic_vector(to_signed(805,16));
ROM(591) <= std_logic_vector(to_signed(806,16));
ROM(592) <= std_logic_vector(to_signed(807,16));
ROM(593) <= std_logic_vector(to_signed(808,16));
ROM(594) <= std_logic_vector(to_signed(809,16));
ROM(595) <= std_logic_vector(to_signed(810,16));
ROM(596) <= std_logic_vector(to_signed(811,16));
ROM(597) <= std_logic_vector(to_signed(812,16));
ROM(598) <= std_logic_vector(to_signed(813,16));
ROM(599) <= std_logic_vector(to_signed(814,16));
ROM(600) <= std_logic_vector(to_signed(815,16));
ROM(601) <= std_logic_vector(to_signed(816,16));
ROM(602) <= std_logic_vector(to_signed(817,16));
ROM(603) <= std_logic_vector(to_signed(818,16));
ROM(604) <= std_logic_vector(to_signed(819,16));
ROM(605) <= std_logic_vector(to_signed(820,16));
ROM(606) <= std_logic_vector(to_signed(821,16));
ROM(607) <= std_logic_vector(to_signed(822,16));
ROM(608) <= std_logic_vector(to_signed(822,16));
ROM(609) <= std_logic_vector(to_signed(823,16));
ROM(610) <= std_logic_vector(to_signed(824,16));
ROM(611) <= std_logic_vector(to_signed(825,16));
ROM(612) <= std_logic_vector(to_signed(826,16));
ROM(613) <= std_logic_vector(to_signed(827,16));
ROM(614) <= std_logic_vector(to_signed(828,16));
ROM(615) <= std_logic_vector(to_signed(829,16));
ROM(616) <= std_logic_vector(to_signed(830,16));
ROM(617) <= std_logic_vector(to_signed(831,16));
ROM(618) <= std_logic_vector(to_signed(832,16));
ROM(619) <= std_logic_vector(to_signed(833,16));
ROM(620) <= std_logic_vector(to_signed(834,16));
ROM(621) <= std_logic_vector(to_signed(834,16));
ROM(622) <= std_logic_vector(to_signed(835,16));
ROM(623) <= std_logic_vector(to_signed(836,16));
ROM(624) <= std_logic_vector(to_signed(837,16));
ROM(625) <= std_logic_vector(to_signed(838,16));
ROM(626) <= std_logic_vector(to_signed(839,16));
ROM(627) <= std_logic_vector(to_signed(840,16));
ROM(628) <= std_logic_vector(to_signed(841,16));
ROM(629) <= std_logic_vector(to_signed(842,16));
ROM(630) <= std_logic_vector(to_signed(843,16));
ROM(631) <= std_logic_vector(to_signed(843,16));
ROM(632) <= std_logic_vector(to_signed(844,16));
ROM(633) <= std_logic_vector(to_signed(845,16));
ROM(634) <= std_logic_vector(to_signed(846,16));
ROM(635) <= std_logic_vector(to_signed(847,16));
ROM(636) <= std_logic_vector(to_signed(848,16));
ROM(637) <= std_logic_vector(to_signed(849,16));
ROM(638) <= std_logic_vector(to_signed(850,16));
ROM(639) <= std_logic_vector(to_signed(851,16));
ROM(640) <= std_logic_vector(to_signed(851,16));
ROM(641) <= std_logic_vector(to_signed(852,16));
ROM(642) <= std_logic_vector(to_signed(853,16));
ROM(643) <= std_logic_vector(to_signed(854,16));
ROM(644) <= std_logic_vector(to_signed(855,16));
ROM(645) <= std_logic_vector(to_signed(856,16));
ROM(646) <= std_logic_vector(to_signed(857,16));
ROM(647) <= std_logic_vector(to_signed(857,16));
ROM(648) <= std_logic_vector(to_signed(858,16));
ROM(649) <= std_logic_vector(to_signed(859,16));
ROM(650) <= std_logic_vector(to_signed(860,16));
ROM(651) <= std_logic_vector(to_signed(861,16));
ROM(652) <= std_logic_vector(to_signed(862,16));
ROM(653) <= std_logic_vector(to_signed(863,16));
ROM(654) <= std_logic_vector(to_signed(863,16));
ROM(655) <= std_logic_vector(to_signed(864,16));
ROM(656) <= std_logic_vector(to_signed(865,16));
ROM(657) <= std_logic_vector(to_signed(866,16));
ROM(658) <= std_logic_vector(to_signed(867,16));
ROM(659) <= std_logic_vector(to_signed(868,16));
ROM(660) <= std_logic_vector(to_signed(868,16));
ROM(661) <= std_logic_vector(to_signed(869,16));
ROM(662) <= std_logic_vector(to_signed(870,16));
ROM(663) <= std_logic_vector(to_signed(871,16));
ROM(664) <= std_logic_vector(to_signed(872,16));
ROM(665) <= std_logic_vector(to_signed(873,16));
ROM(666) <= std_logic_vector(to_signed(873,16));
ROM(667) <= std_logic_vector(to_signed(874,16));
ROM(668) <= std_logic_vector(to_signed(875,16));
ROM(669) <= std_logic_vector(to_signed(876,16));
ROM(670) <= std_logic_vector(to_signed(877,16));
ROM(671) <= std_logic_vector(to_signed(878,16));
ROM(672) <= std_logic_vector(to_signed(878,16));
ROM(673) <= std_logic_vector(to_signed(879,16));
ROM(674) <= std_logic_vector(to_signed(880,16));
ROM(675) <= std_logic_vector(to_signed(881,16));
ROM(676) <= std_logic_vector(to_signed(882,16));
ROM(677) <= std_logic_vector(to_signed(882,16));
ROM(678) <= std_logic_vector(to_signed(883,16));
ROM(679) <= std_logic_vector(to_signed(884,16));
ROM(680) <= std_logic_vector(to_signed(885,16));
ROM(681) <= std_logic_vector(to_signed(885,16));
ROM(682) <= std_logic_vector(to_signed(886,16));
ROM(683) <= std_logic_vector(to_signed(887,16));
ROM(684) <= std_logic_vector(to_signed(888,16));
ROM(685) <= std_logic_vector(to_signed(889,16));
ROM(686) <= std_logic_vector(to_signed(889,16));
ROM(687) <= std_logic_vector(to_signed(890,16));
ROM(688) <= std_logic_vector(to_signed(891,16));
ROM(689) <= std_logic_vector(to_signed(892,16));
ROM(690) <= std_logic_vector(to_signed(893,16));
ROM(691) <= std_logic_vector(to_signed(893,16));
ROM(692) <= std_logic_vector(to_signed(894,16));
ROM(693) <= std_logic_vector(to_signed(895,16));
ROM(694) <= std_logic_vector(to_signed(896,16));
ROM(695) <= std_logic_vector(to_signed(896,16));
ROM(696) <= std_logic_vector(to_signed(897,16));
ROM(697) <= std_logic_vector(to_signed(898,16));
ROM(698) <= std_logic_vector(to_signed(899,16));
ROM(699) <= std_logic_vector(to_signed(899,16));
ROM(700) <= std_logic_vector(to_signed(900,16));
ROM(701) <= std_logic_vector(to_signed(901,16));
ROM(702) <= std_logic_vector(to_signed(902,16));
ROM(703) <= std_logic_vector(to_signed(902,16));
ROM(704) <= std_logic_vector(to_signed(903,16));
ROM(705) <= std_logic_vector(to_signed(904,16));
ROM(706) <= std_logic_vector(to_signed(905,16));
ROM(707) <= std_logic_vector(to_signed(905,16));
ROM(708) <= std_logic_vector(to_signed(906,16));
ROM(709) <= std_logic_vector(to_signed(907,16));
ROM(710) <= std_logic_vector(to_signed(907,16));
ROM(711) <= std_logic_vector(to_signed(908,16));
ROM(712) <= std_logic_vector(to_signed(909,16));
ROM(713) <= std_logic_vector(to_signed(910,16));
ROM(714) <= std_logic_vector(to_signed(910,16));
ROM(715) <= std_logic_vector(to_signed(911,16));
ROM(716) <= std_logic_vector(to_signed(912,16));
ROM(717) <= std_logic_vector(to_signed(913,16));
ROM(718) <= std_logic_vector(to_signed(913,16));
ROM(719) <= std_logic_vector(to_signed(914,16));
ROM(720) <= std_logic_vector(to_signed(915,16));
ROM(721) <= std_logic_vector(to_signed(915,16));
ROM(722) <= std_logic_vector(to_signed(916,16));
ROM(723) <= std_logic_vector(to_signed(917,16));
ROM(724) <= std_logic_vector(to_signed(917,16));
ROM(725) <= std_logic_vector(to_signed(918,16));
ROM(726) <= std_logic_vector(to_signed(919,16));
ROM(727) <= std_logic_vector(to_signed(920,16));
ROM(728) <= std_logic_vector(to_signed(920,16));
ROM(729) <= std_logic_vector(to_signed(921,16));
ROM(730) <= std_logic_vector(to_signed(922,16));
ROM(731) <= std_logic_vector(to_signed(922,16));
ROM(732) <= std_logic_vector(to_signed(923,16));
ROM(733) <= std_logic_vector(to_signed(924,16));
ROM(734) <= std_logic_vector(to_signed(924,16));
ROM(735) <= std_logic_vector(to_signed(925,16));
ROM(736) <= std_logic_vector(to_signed(926,16));
ROM(737) <= std_logic_vector(to_signed(926,16));
ROM(738) <= std_logic_vector(to_signed(927,16));
ROM(739) <= std_logic_vector(to_signed(928,16));
ROM(740) <= std_logic_vector(to_signed(928,16));
ROM(741) <= std_logic_vector(to_signed(929,16));
ROM(742) <= std_logic_vector(to_signed(930,16));
ROM(743) <= std_logic_vector(to_signed(930,16));
ROM(744) <= std_logic_vector(to_signed(931,16));
ROM(745) <= std_logic_vector(to_signed(932,16));
ROM(746) <= std_logic_vector(to_signed(932,16));
ROM(747) <= std_logic_vector(to_signed(933,16));
ROM(748) <= std_logic_vector(to_signed(934,16));
ROM(749) <= std_logic_vector(to_signed(934,16));
ROM(750) <= std_logic_vector(to_signed(935,16));
ROM(751) <= std_logic_vector(to_signed(936,16));
ROM(752) <= std_logic_vector(to_signed(936,16));
ROM(753) <= std_logic_vector(to_signed(937,16));
ROM(754) <= std_logic_vector(to_signed(937,16));
ROM(755) <= std_logic_vector(to_signed(938,16));
ROM(756) <= std_logic_vector(to_signed(939,16));
ROM(757) <= std_logic_vector(to_signed(939,16));
ROM(758) <= std_logic_vector(to_signed(940,16));
ROM(759) <= std_logic_vector(to_signed(941,16));
ROM(760) <= std_logic_vector(to_signed(941,16));
ROM(761) <= std_logic_vector(to_signed(942,16));
ROM(762) <= std_logic_vector(to_signed(942,16));
ROM(763) <= std_logic_vector(to_signed(943,16));
ROM(764) <= std_logic_vector(to_signed(944,16));
ROM(765) <= std_logic_vector(to_signed(944,16));
ROM(766) <= std_logic_vector(to_signed(945,16));
ROM(767) <= std_logic_vector(to_signed(945,16));
ROM(768) <= std_logic_vector(to_signed(946,16));
ROM(769) <= std_logic_vector(to_signed(947,16));
ROM(770) <= std_logic_vector(to_signed(947,16));
ROM(771) <= std_logic_vector(to_signed(948,16));
ROM(772) <= std_logic_vector(to_signed(948,16));
ROM(773) <= std_logic_vector(to_signed(949,16));
ROM(774) <= std_logic_vector(to_signed(950,16));
ROM(775) <= std_logic_vector(to_signed(950,16));
ROM(776) <= std_logic_vector(to_signed(951,16));
ROM(777) <= std_logic_vector(to_signed(951,16));
ROM(778) <= std_logic_vector(to_signed(952,16));
ROM(779) <= std_logic_vector(to_signed(953,16));
ROM(780) <= std_logic_vector(to_signed(953,16));
ROM(781) <= std_logic_vector(to_signed(954,16));
ROM(782) <= std_logic_vector(to_signed(954,16));
ROM(783) <= std_logic_vector(to_signed(955,16));
ROM(784) <= std_logic_vector(to_signed(955,16));
ROM(785) <= std_logic_vector(to_signed(956,16));
ROM(786) <= std_logic_vector(to_signed(957,16));
ROM(787) <= std_logic_vector(to_signed(957,16));
ROM(788) <= std_logic_vector(to_signed(958,16));
ROM(789) <= std_logic_vector(to_signed(958,16));
ROM(790) <= std_logic_vector(to_signed(959,16));
ROM(791) <= std_logic_vector(to_signed(959,16));
ROM(792) <= std_logic_vector(to_signed(960,16));
ROM(793) <= std_logic_vector(to_signed(960,16));
ROM(794) <= std_logic_vector(to_signed(961,16));
ROM(795) <= std_logic_vector(to_signed(961,16));
ROM(796) <= std_logic_vector(to_signed(962,16));
ROM(797) <= std_logic_vector(to_signed(963,16));
ROM(798) <= std_logic_vector(to_signed(963,16));
ROM(799) <= std_logic_vector(to_signed(964,16));
ROM(800) <= std_logic_vector(to_signed(964,16));
ROM(801) <= std_logic_vector(to_signed(965,16));
ROM(802) <= std_logic_vector(to_signed(965,16));
ROM(803) <= std_logic_vector(to_signed(966,16));
ROM(804) <= std_logic_vector(to_signed(966,16));
ROM(805) <= std_logic_vector(to_signed(967,16));
ROM(806) <= std_logic_vector(to_signed(967,16));
ROM(807) <= std_logic_vector(to_signed(968,16));
ROM(808) <= std_logic_vector(to_signed(968,16));
ROM(809) <= std_logic_vector(to_signed(969,16));
ROM(810) <= std_logic_vector(to_signed(969,16));
ROM(811) <= std_logic_vector(to_signed(970,16));
ROM(812) <= std_logic_vector(to_signed(970,16));
ROM(813) <= std_logic_vector(to_signed(971,16));
ROM(814) <= std_logic_vector(to_signed(971,16));
ROM(815) <= std_logic_vector(to_signed(972,16));
ROM(816) <= std_logic_vector(to_signed(972,16));
ROM(817) <= std_logic_vector(to_signed(973,16));
ROM(818) <= std_logic_vector(to_signed(973,16));
ROM(819) <= std_logic_vector(to_signed(974,16));
ROM(820) <= std_logic_vector(to_signed(974,16));
ROM(821) <= std_logic_vector(to_signed(975,16));
ROM(822) <= std_logic_vector(to_signed(975,16));
ROM(823) <= std_logic_vector(to_signed(976,16));
ROM(824) <= std_logic_vector(to_signed(976,16));
ROM(825) <= std_logic_vector(to_signed(977,16));
ROM(826) <= std_logic_vector(to_signed(977,16));
ROM(827) <= std_logic_vector(to_signed(978,16));
ROM(828) <= std_logic_vector(to_signed(978,16));
ROM(829) <= std_logic_vector(to_signed(979,16));
ROM(830) <= std_logic_vector(to_signed(979,16));
ROM(831) <= std_logic_vector(to_signed(979,16));
ROM(832) <= std_logic_vector(to_signed(980,16));
ROM(833) <= std_logic_vector(to_signed(980,16));
ROM(834) <= std_logic_vector(to_signed(981,16));
ROM(835) <= std_logic_vector(to_signed(981,16));
ROM(836) <= std_logic_vector(to_signed(982,16));
ROM(837) <= std_logic_vector(to_signed(982,16));
ROM(838) <= std_logic_vector(to_signed(983,16));
ROM(839) <= std_logic_vector(to_signed(983,16));
ROM(840) <= std_logic_vector(to_signed(983,16));
ROM(841) <= std_logic_vector(to_signed(984,16));
ROM(842) <= std_logic_vector(to_signed(984,16));
ROM(843) <= std_logic_vector(to_signed(985,16));
ROM(844) <= std_logic_vector(to_signed(985,16));
ROM(845) <= std_logic_vector(to_signed(986,16));
ROM(846) <= std_logic_vector(to_signed(986,16));
ROM(847) <= std_logic_vector(to_signed(986,16));
ROM(848) <= std_logic_vector(to_signed(987,16));
ROM(849) <= std_logic_vector(to_signed(987,16));
ROM(850) <= std_logic_vector(to_signed(988,16));
ROM(851) <= std_logic_vector(to_signed(988,16));
ROM(852) <= std_logic_vector(to_signed(989,16));
ROM(853) <= std_logic_vector(to_signed(989,16));
ROM(854) <= std_logic_vector(to_signed(989,16));
ROM(855) <= std_logic_vector(to_signed(990,16));
ROM(856) <= std_logic_vector(to_signed(990,16));
ROM(857) <= std_logic_vector(to_signed(991,16));
ROM(858) <= std_logic_vector(to_signed(991,16));
ROM(859) <= std_logic_vector(to_signed(991,16));
ROM(860) <= std_logic_vector(to_signed(992,16));
ROM(861) <= std_logic_vector(to_signed(992,16));
ROM(862) <= std_logic_vector(to_signed(993,16));
ROM(863) <= std_logic_vector(to_signed(993,16));
ROM(864) <= std_logic_vector(to_signed(993,16));
ROM(865) <= std_logic_vector(to_signed(994,16));
ROM(866) <= std_logic_vector(to_signed(994,16));
ROM(867) <= std_logic_vector(to_signed(994,16));
ROM(868) <= std_logic_vector(to_signed(995,16));
ROM(869) <= std_logic_vector(to_signed(995,16));
ROM(870) <= std_logic_vector(to_signed(996,16));
ROM(871) <= std_logic_vector(to_signed(996,16));
ROM(872) <= std_logic_vector(to_signed(996,16));
ROM(873) <= std_logic_vector(to_signed(997,16));
ROM(874) <= std_logic_vector(to_signed(997,16));
ROM(875) <= std_logic_vector(to_signed(997,16));
ROM(876) <= std_logic_vector(to_signed(998,16));
ROM(877) <= std_logic_vector(to_signed(998,16));
ROM(878) <= std_logic_vector(to_signed(998,16));
ROM(879) <= std_logic_vector(to_signed(999,16));
ROM(880) <= std_logic_vector(to_signed(999,16));
ROM(881) <= std_logic_vector(to_signed(999,16));
ROM(882) <= std_logic_vector(to_signed(1000,16));
ROM(883) <= std_logic_vector(to_signed(1000,16));
ROM(884) <= std_logic_vector(to_signed(1000,16));
ROM(885) <= std_logic_vector(to_signed(1001,16));
ROM(886) <= std_logic_vector(to_signed(1001,16));
ROM(887) <= std_logic_vector(to_signed(1001,16));
ROM(888) <= std_logic_vector(to_signed(1002,16));
ROM(889) <= std_logic_vector(to_signed(1002,16));
ROM(890) <= std_logic_vector(to_signed(1002,16));
ROM(891) <= std_logic_vector(to_signed(1003,16));
ROM(892) <= std_logic_vector(to_signed(1003,16));
ROM(893) <= std_logic_vector(to_signed(1003,16));
ROM(894) <= std_logic_vector(to_signed(1004,16));
ROM(895) <= std_logic_vector(to_signed(1004,16));
ROM(896) <= std_logic_vector(to_signed(1004,16));
ROM(897) <= std_logic_vector(to_signed(1005,16));
ROM(898) <= std_logic_vector(to_signed(1005,16));
ROM(899) <= std_logic_vector(to_signed(1005,16));
ROM(900) <= std_logic_vector(to_signed(1006,16));
ROM(901) <= std_logic_vector(to_signed(1006,16));
ROM(902) <= std_logic_vector(to_signed(1006,16));
ROM(903) <= std_logic_vector(to_signed(1006,16));
ROM(904) <= std_logic_vector(to_signed(1007,16));
ROM(905) <= std_logic_vector(to_signed(1007,16));
ROM(906) <= std_logic_vector(to_signed(1007,16));
ROM(907) <= std_logic_vector(to_signed(1008,16));
ROM(908) <= std_logic_vector(to_signed(1008,16));
ROM(909) <= std_logic_vector(to_signed(1008,16));
ROM(910) <= std_logic_vector(to_signed(1008,16));
ROM(911) <= std_logic_vector(to_signed(1009,16));
ROM(912) <= std_logic_vector(to_signed(1009,16));
ROM(913) <= std_logic_vector(to_signed(1009,16));
ROM(914) <= std_logic_vector(to_signed(1009,16));
ROM(915) <= std_logic_vector(to_signed(1010,16));
ROM(916) <= std_logic_vector(to_signed(1010,16));
ROM(917) <= std_logic_vector(to_signed(1010,16));
ROM(918) <= std_logic_vector(to_signed(1010,16));
ROM(919) <= std_logic_vector(to_signed(1011,16));
ROM(920) <= std_logic_vector(to_signed(1011,16));
ROM(921) <= std_logic_vector(to_signed(1011,16));
ROM(922) <= std_logic_vector(to_signed(1011,16));
ROM(923) <= std_logic_vector(to_signed(1012,16));
ROM(924) <= std_logic_vector(to_signed(1012,16));
ROM(925) <= std_logic_vector(to_signed(1012,16));
ROM(926) <= std_logic_vector(to_signed(1012,16));
ROM(927) <= std_logic_vector(to_signed(1013,16));
ROM(928) <= std_logic_vector(to_signed(1013,16));
ROM(929) <= std_logic_vector(to_signed(1013,16));
ROM(930) <= std_logic_vector(to_signed(1013,16));
ROM(931) <= std_logic_vector(to_signed(1014,16));
ROM(932) <= std_logic_vector(to_signed(1014,16));
ROM(933) <= std_logic_vector(to_signed(1014,16));
ROM(934) <= std_logic_vector(to_signed(1014,16));
ROM(935) <= std_logic_vector(to_signed(1014,16));
ROM(936) <= std_logic_vector(to_signed(1015,16));
ROM(937) <= std_logic_vector(to_signed(1015,16));
ROM(938) <= std_logic_vector(to_signed(1015,16));
ROM(939) <= std_logic_vector(to_signed(1015,16));
ROM(940) <= std_logic_vector(to_signed(1016,16));
ROM(941) <= std_logic_vector(to_signed(1016,16));
ROM(942) <= std_logic_vector(to_signed(1016,16));
ROM(943) <= std_logic_vector(to_signed(1016,16));
ROM(944) <= std_logic_vector(to_signed(1016,16));
ROM(945) <= std_logic_vector(to_signed(1016,16));
ROM(946) <= std_logic_vector(to_signed(1017,16));
ROM(947) <= std_logic_vector(to_signed(1017,16));
ROM(948) <= std_logic_vector(to_signed(1017,16));
ROM(949) <= std_logic_vector(to_signed(1017,16));
ROM(950) <= std_logic_vector(to_signed(1017,16));
ROM(951) <= std_logic_vector(to_signed(1018,16));
ROM(952) <= std_logic_vector(to_signed(1018,16));
ROM(953) <= std_logic_vector(to_signed(1018,16));
ROM(954) <= std_logic_vector(to_signed(1018,16));
ROM(955) <= std_logic_vector(to_signed(1018,16));
ROM(956) <= std_logic_vector(to_signed(1018,16));
ROM(957) <= std_logic_vector(to_signed(1019,16));
ROM(958) <= std_logic_vector(to_signed(1019,16));
ROM(959) <= std_logic_vector(to_signed(1019,16));
ROM(960) <= std_logic_vector(to_signed(1019,16));
ROM(961) <= std_logic_vector(to_signed(1019,16));
ROM(962) <= std_logic_vector(to_signed(1019,16));
ROM(963) <= std_logic_vector(to_signed(1020,16));
ROM(964) <= std_logic_vector(to_signed(1020,16));
ROM(965) <= std_logic_vector(to_signed(1020,16));
ROM(966) <= std_logic_vector(to_signed(1020,16));
ROM(967) <= std_logic_vector(to_signed(1020,16));
ROM(968) <= std_logic_vector(to_signed(1020,16));
ROM(969) <= std_logic_vector(to_signed(1020,16));
ROM(970) <= std_logic_vector(to_signed(1020,16));
ROM(971) <= std_logic_vector(to_signed(1021,16));
ROM(972) <= std_logic_vector(to_signed(1021,16));
ROM(973) <= std_logic_vector(to_signed(1021,16));
ROM(974) <= std_logic_vector(to_signed(1021,16));
ROM(975) <= std_logic_vector(to_signed(1021,16));
ROM(976) <= std_logic_vector(to_signed(1021,16));
ROM(977) <= std_logic_vector(to_signed(1021,16));
ROM(978) <= std_logic_vector(to_signed(1021,16));
ROM(979) <= std_logic_vector(to_signed(1022,16));
ROM(980) <= std_logic_vector(to_signed(1022,16));
ROM(981) <= std_logic_vector(to_signed(1022,16));
ROM(982) <= std_logic_vector(to_signed(1022,16));
ROM(983) <= std_logic_vector(to_signed(1022,16));
ROM(984) <= std_logic_vector(to_signed(1022,16));
ROM(985) <= std_logic_vector(to_signed(1022,16));
ROM(986) <= std_logic_vector(to_signed(1022,16));
ROM(987) <= std_logic_vector(to_signed(1022,16));
ROM(988) <= std_logic_vector(to_signed(1022,16));
ROM(989) <= std_logic_vector(to_signed(1023,16));
ROM(990) <= std_logic_vector(to_signed(1023,16));
ROM(991) <= std_logic_vector(to_signed(1023,16));
ROM(992) <= std_logic_vector(to_signed(1023,16));
ROM(993) <= std_logic_vector(to_signed(1023,16));
ROM(994) <= std_logic_vector(to_signed(1023,16));
ROM(995) <= std_logic_vector(to_signed(1023,16));
ROM(996) <= std_logic_vector(to_signed(1023,16));
ROM(997) <= std_logic_vector(to_signed(1023,16));
ROM(998) <= std_logic_vector(to_signed(1023,16));
ROM(999) <= std_logic_vector(to_signed(1023,16));
ROM(1000) <= std_logic_vector(to_signed(1023,16));
ROM(1001) <= std_logic_vector(to_signed(1023,16));
ROM(1002) <= std_logic_vector(to_signed(1023,16));
ROM(1003) <= std_logic_vector(to_signed(1023,16));
ROM(1004) <= std_logic_vector(to_signed(1024,16));
ROM(1005) <= std_logic_vector(to_signed(1024,16));
ROM(1006) <= std_logic_vector(to_signed(1024,16));
ROM(1007) <= std_logic_vector(to_signed(1024,16));
ROM(1008) <= std_logic_vector(to_signed(1024,16));
ROM(1009) <= std_logic_vector(to_signed(1024,16));
ROM(1010) <= std_logic_vector(to_signed(1024,16));
ROM(1011) <= std_logic_vector(to_signed(1024,16));
ROM(1012) <= std_logic_vector(to_signed(1024,16));
ROM(1013) <= std_logic_vector(to_signed(1024,16));
ROM(1014) <= std_logic_vector(to_signed(1024,16));
ROM(1015) <= std_logic_vector(to_signed(1024,16));
ROM(1016) <= std_logic_vector(to_signed(1024,16));
ROM(1017) <= std_logic_vector(to_signed(1024,16));
ROM(1018) <= std_logic_vector(to_signed(1024,16));
ROM(1019) <= std_logic_vector(to_signed(1024,16));
ROM(1020) <= std_logic_vector(to_signed(1024,16));
ROM(1021) <= std_logic_vector(to_signed(1024,16));
ROM(1022) <= std_logic_vector(to_signed(1024,16));
ROM(1023) <= std_logic_vector(to_signed(1024,16));
ROM(1024) <= std_logic_vector(to_signed(1024,16));
ROM(1025) <= std_logic_vector(to_signed(1024,16));
ROM(1026) <= std_logic_vector(to_signed(1024,16));
ROM(1027) <= std_logic_vector(to_signed(1024,16));
ROM(1028) <= std_logic_vector(to_signed(1024,16));
ROM(1029) <= std_logic_vector(to_signed(1024,16));
ROM(1030) <= std_logic_vector(to_signed(1024,16));
ROM(1031) <= std_logic_vector(to_signed(1024,16));
ROM(1032) <= std_logic_vector(to_signed(1024,16));
ROM(1033) <= std_logic_vector(to_signed(1024,16));
ROM(1034) <= std_logic_vector(to_signed(1024,16));
ROM(1035) <= std_logic_vector(to_signed(1024,16));
ROM(1036) <= std_logic_vector(to_signed(1024,16));
ROM(1037) <= std_logic_vector(to_signed(1024,16));
ROM(1038) <= std_logic_vector(to_signed(1024,16));
ROM(1039) <= std_logic_vector(to_signed(1024,16));
ROM(1040) <= std_logic_vector(to_signed(1024,16));
ROM(1041) <= std_logic_vector(to_signed(1024,16));
ROM(1042) <= std_logic_vector(to_signed(1024,16));
ROM(1043) <= std_logic_vector(to_signed(1024,16));
ROM(1044) <= std_logic_vector(to_signed(1024,16));
ROM(1045) <= std_logic_vector(to_signed(1023,16));
ROM(1046) <= std_logic_vector(to_signed(1023,16));
ROM(1047) <= std_logic_vector(to_signed(1023,16));
ROM(1048) <= std_logic_vector(to_signed(1023,16));
ROM(1049) <= std_logic_vector(to_signed(1023,16));
ROM(1050) <= std_logic_vector(to_signed(1023,16));
ROM(1051) <= std_logic_vector(to_signed(1023,16));
ROM(1052) <= std_logic_vector(to_signed(1023,16));
ROM(1053) <= std_logic_vector(to_signed(1023,16));
ROM(1054) <= std_logic_vector(to_signed(1023,16));
ROM(1055) <= std_logic_vector(to_signed(1023,16));
ROM(1056) <= std_logic_vector(to_signed(1023,16));
ROM(1057) <= std_logic_vector(to_signed(1023,16));
ROM(1058) <= std_logic_vector(to_signed(1023,16));
ROM(1059) <= std_logic_vector(to_signed(1023,16));
ROM(1060) <= std_logic_vector(to_signed(1022,16));
ROM(1061) <= std_logic_vector(to_signed(1022,16));
ROM(1062) <= std_logic_vector(to_signed(1022,16));
ROM(1063) <= std_logic_vector(to_signed(1022,16));
ROM(1064) <= std_logic_vector(to_signed(1022,16));
ROM(1065) <= std_logic_vector(to_signed(1022,16));
ROM(1066) <= std_logic_vector(to_signed(1022,16));
ROM(1067) <= std_logic_vector(to_signed(1022,16));
ROM(1068) <= std_logic_vector(to_signed(1022,16));
ROM(1069) <= std_logic_vector(to_signed(1022,16));
ROM(1070) <= std_logic_vector(to_signed(1021,16));
ROM(1071) <= std_logic_vector(to_signed(1021,16));
ROM(1072) <= std_logic_vector(to_signed(1021,16));
ROM(1073) <= std_logic_vector(to_signed(1021,16));
ROM(1074) <= std_logic_vector(to_signed(1021,16));
ROM(1075) <= std_logic_vector(to_signed(1021,16));
ROM(1076) <= std_logic_vector(to_signed(1021,16));
ROM(1077) <= std_logic_vector(to_signed(1021,16));
ROM(1078) <= std_logic_vector(to_signed(1020,16));
ROM(1079) <= std_logic_vector(to_signed(1020,16));
ROM(1080) <= std_logic_vector(to_signed(1020,16));
ROM(1081) <= std_logic_vector(to_signed(1020,16));
ROM(1082) <= std_logic_vector(to_signed(1020,16));
ROM(1083) <= std_logic_vector(to_signed(1020,16));
ROM(1084) <= std_logic_vector(to_signed(1020,16));
ROM(1085) <= std_logic_vector(to_signed(1020,16));
ROM(1086) <= std_logic_vector(to_signed(1019,16));
ROM(1087) <= std_logic_vector(to_signed(1019,16));
ROM(1088) <= std_logic_vector(to_signed(1019,16));
ROM(1089) <= std_logic_vector(to_signed(1019,16));
ROM(1090) <= std_logic_vector(to_signed(1019,16));
ROM(1091) <= std_logic_vector(to_signed(1019,16));
ROM(1092) <= std_logic_vector(to_signed(1018,16));
ROM(1093) <= std_logic_vector(to_signed(1018,16));
ROM(1094) <= std_logic_vector(to_signed(1018,16));
ROM(1095) <= std_logic_vector(to_signed(1018,16));
ROM(1096) <= std_logic_vector(to_signed(1018,16));
ROM(1097) <= std_logic_vector(to_signed(1018,16));
ROM(1098) <= std_logic_vector(to_signed(1017,16));
ROM(1099) <= std_logic_vector(to_signed(1017,16));
ROM(1100) <= std_logic_vector(to_signed(1017,16));
ROM(1101) <= std_logic_vector(to_signed(1017,16));
ROM(1102) <= std_logic_vector(to_signed(1017,16));
ROM(1103) <= std_logic_vector(to_signed(1016,16));
ROM(1104) <= std_logic_vector(to_signed(1016,16));
ROM(1105) <= std_logic_vector(to_signed(1016,16));
ROM(1106) <= std_logic_vector(to_signed(1016,16));
ROM(1107) <= std_logic_vector(to_signed(1016,16));
ROM(1108) <= std_logic_vector(to_signed(1016,16));
ROM(1109) <= std_logic_vector(to_signed(1015,16));
ROM(1110) <= std_logic_vector(to_signed(1015,16));
ROM(1111) <= std_logic_vector(to_signed(1015,16));
ROM(1112) <= std_logic_vector(to_signed(1015,16));
ROM(1113) <= std_logic_vector(to_signed(1014,16));
ROM(1114) <= std_logic_vector(to_signed(1014,16));
ROM(1115) <= std_logic_vector(to_signed(1014,16));
ROM(1116) <= std_logic_vector(to_signed(1014,16));
ROM(1117) <= std_logic_vector(to_signed(1014,16));
ROM(1118) <= std_logic_vector(to_signed(1013,16));
ROM(1119) <= std_logic_vector(to_signed(1013,16));
ROM(1120) <= std_logic_vector(to_signed(1013,16));
ROM(1121) <= std_logic_vector(to_signed(1013,16));
ROM(1122) <= std_logic_vector(to_signed(1012,16));
ROM(1123) <= std_logic_vector(to_signed(1012,16));
ROM(1124) <= std_logic_vector(to_signed(1012,16));
ROM(1125) <= std_logic_vector(to_signed(1012,16));
ROM(1126) <= std_logic_vector(to_signed(1011,16));
ROM(1127) <= std_logic_vector(to_signed(1011,16));
ROM(1128) <= std_logic_vector(to_signed(1011,16));
ROM(1129) <= std_logic_vector(to_signed(1011,16));
ROM(1130) <= std_logic_vector(to_signed(1010,16));
ROM(1131) <= std_logic_vector(to_signed(1010,16));
ROM(1132) <= std_logic_vector(to_signed(1010,16));
ROM(1133) <= std_logic_vector(to_signed(1010,16));
ROM(1134) <= std_logic_vector(to_signed(1009,16));
ROM(1135) <= std_logic_vector(to_signed(1009,16));
ROM(1136) <= std_logic_vector(to_signed(1009,16));
ROM(1137) <= std_logic_vector(to_signed(1009,16));
ROM(1138) <= std_logic_vector(to_signed(1008,16));
ROM(1139) <= std_logic_vector(to_signed(1008,16));
ROM(1140) <= std_logic_vector(to_signed(1008,16));
ROM(1141) <= std_logic_vector(to_signed(1008,16));
ROM(1142) <= std_logic_vector(to_signed(1007,16));
ROM(1143) <= std_logic_vector(to_signed(1007,16));
ROM(1144) <= std_logic_vector(to_signed(1007,16));
ROM(1145) <= std_logic_vector(to_signed(1006,16));
ROM(1146) <= std_logic_vector(to_signed(1006,16));
ROM(1147) <= std_logic_vector(to_signed(1006,16));
ROM(1148) <= std_logic_vector(to_signed(1006,16));
ROM(1149) <= std_logic_vector(to_signed(1005,16));
ROM(1150) <= std_logic_vector(to_signed(1005,16));
ROM(1151) <= std_logic_vector(to_signed(1005,16));
ROM(1152) <= std_logic_vector(to_signed(1004,16));
ROM(1153) <= std_logic_vector(to_signed(1004,16));
ROM(1154) <= std_logic_vector(to_signed(1004,16));
ROM(1155) <= std_logic_vector(to_signed(1003,16));
ROM(1156) <= std_logic_vector(to_signed(1003,16));
ROM(1157) <= std_logic_vector(to_signed(1003,16));
ROM(1158) <= std_logic_vector(to_signed(1002,16));
ROM(1159) <= std_logic_vector(to_signed(1002,16));
ROM(1160) <= std_logic_vector(to_signed(1002,16));
ROM(1161) <= std_logic_vector(to_signed(1001,16));
ROM(1162) <= std_logic_vector(to_signed(1001,16));
ROM(1163) <= std_logic_vector(to_signed(1001,16));
ROM(1164) <= std_logic_vector(to_signed(1000,16));
ROM(1165) <= std_logic_vector(to_signed(1000,16));
ROM(1166) <= std_logic_vector(to_signed(1000,16));
ROM(1167) <= std_logic_vector(to_signed(999,16));
ROM(1168) <= std_logic_vector(to_signed(999,16));
ROM(1169) <= std_logic_vector(to_signed(999,16));
ROM(1170) <= std_logic_vector(to_signed(998,16));
ROM(1171) <= std_logic_vector(to_signed(998,16));
ROM(1172) <= std_logic_vector(to_signed(998,16));
ROM(1173) <= std_logic_vector(to_signed(997,16));
ROM(1174) <= std_logic_vector(to_signed(997,16));
ROM(1175) <= std_logic_vector(to_signed(997,16));
ROM(1176) <= std_logic_vector(to_signed(996,16));
ROM(1177) <= std_logic_vector(to_signed(996,16));
ROM(1178) <= std_logic_vector(to_signed(996,16));
ROM(1179) <= std_logic_vector(to_signed(995,16));
ROM(1180) <= std_logic_vector(to_signed(995,16));
ROM(1181) <= std_logic_vector(to_signed(994,16));
ROM(1182) <= std_logic_vector(to_signed(994,16));
ROM(1183) <= std_logic_vector(to_signed(994,16));
ROM(1184) <= std_logic_vector(to_signed(993,16));
ROM(1185) <= std_logic_vector(to_signed(993,16));
ROM(1186) <= std_logic_vector(to_signed(993,16));
ROM(1187) <= std_logic_vector(to_signed(992,16));
ROM(1188) <= std_logic_vector(to_signed(992,16));
ROM(1189) <= std_logic_vector(to_signed(991,16));
ROM(1190) <= std_logic_vector(to_signed(991,16));
ROM(1191) <= std_logic_vector(to_signed(991,16));
ROM(1192) <= std_logic_vector(to_signed(990,16));
ROM(1193) <= std_logic_vector(to_signed(990,16));
ROM(1194) <= std_logic_vector(to_signed(989,16));
ROM(1195) <= std_logic_vector(to_signed(989,16));
ROM(1196) <= std_logic_vector(to_signed(989,16));
ROM(1197) <= std_logic_vector(to_signed(988,16));
ROM(1198) <= std_logic_vector(to_signed(988,16));
ROM(1199) <= std_logic_vector(to_signed(987,16));
ROM(1200) <= std_logic_vector(to_signed(987,16));
ROM(1201) <= std_logic_vector(to_signed(986,16));
ROM(1202) <= std_logic_vector(to_signed(986,16));
ROM(1203) <= std_logic_vector(to_signed(986,16));
ROM(1204) <= std_logic_vector(to_signed(985,16));
ROM(1205) <= std_logic_vector(to_signed(985,16));
ROM(1206) <= std_logic_vector(to_signed(984,16));
ROM(1207) <= std_logic_vector(to_signed(984,16));
ROM(1208) <= std_logic_vector(to_signed(983,16));
ROM(1209) <= std_logic_vector(to_signed(983,16));
ROM(1210) <= std_logic_vector(to_signed(983,16));
ROM(1211) <= std_logic_vector(to_signed(982,16));
ROM(1212) <= std_logic_vector(to_signed(982,16));
ROM(1213) <= std_logic_vector(to_signed(981,16));
ROM(1214) <= std_logic_vector(to_signed(981,16));
ROM(1215) <= std_logic_vector(to_signed(980,16));
ROM(1216) <= std_logic_vector(to_signed(980,16));
ROM(1217) <= std_logic_vector(to_signed(979,16));
ROM(1218) <= std_logic_vector(to_signed(979,16));
ROM(1219) <= std_logic_vector(to_signed(979,16));
ROM(1220) <= std_logic_vector(to_signed(978,16));
ROM(1221) <= std_logic_vector(to_signed(978,16));
ROM(1222) <= std_logic_vector(to_signed(977,16));
ROM(1223) <= std_logic_vector(to_signed(977,16));
ROM(1224) <= std_logic_vector(to_signed(976,16));
ROM(1225) <= std_logic_vector(to_signed(976,16));
ROM(1226) <= std_logic_vector(to_signed(975,16));
ROM(1227) <= std_logic_vector(to_signed(975,16));
ROM(1228) <= std_logic_vector(to_signed(974,16));
ROM(1229) <= std_logic_vector(to_signed(974,16));
ROM(1230) <= std_logic_vector(to_signed(973,16));
ROM(1231) <= std_logic_vector(to_signed(973,16));
ROM(1232) <= std_logic_vector(to_signed(972,16));
ROM(1233) <= std_logic_vector(to_signed(972,16));
ROM(1234) <= std_logic_vector(to_signed(971,16));
ROM(1235) <= std_logic_vector(to_signed(971,16));
ROM(1236) <= std_logic_vector(to_signed(970,16));
ROM(1237) <= std_logic_vector(to_signed(970,16));
ROM(1238) <= std_logic_vector(to_signed(969,16));
ROM(1239) <= std_logic_vector(to_signed(969,16));
ROM(1240) <= std_logic_vector(to_signed(968,16));
ROM(1241) <= std_logic_vector(to_signed(968,16));
ROM(1242) <= std_logic_vector(to_signed(967,16));
ROM(1243) <= std_logic_vector(to_signed(967,16));
ROM(1244) <= std_logic_vector(to_signed(966,16));
ROM(1245) <= std_logic_vector(to_signed(966,16));
ROM(1246) <= std_logic_vector(to_signed(965,16));
ROM(1247) <= std_logic_vector(to_signed(965,16));
ROM(1248) <= std_logic_vector(to_signed(964,16));
ROM(1249) <= std_logic_vector(to_signed(964,16));
ROM(1250) <= std_logic_vector(to_signed(963,16));
ROM(1251) <= std_logic_vector(to_signed(963,16));
ROM(1252) <= std_logic_vector(to_signed(962,16));
ROM(1253) <= std_logic_vector(to_signed(961,16));
ROM(1254) <= std_logic_vector(to_signed(961,16));
ROM(1255) <= std_logic_vector(to_signed(960,16));
ROM(1256) <= std_logic_vector(to_signed(960,16));
ROM(1257) <= std_logic_vector(to_signed(959,16));
ROM(1258) <= std_logic_vector(to_signed(959,16));
ROM(1259) <= std_logic_vector(to_signed(958,16));
ROM(1260) <= std_logic_vector(to_signed(958,16));
ROM(1261) <= std_logic_vector(to_signed(957,16));
ROM(1262) <= std_logic_vector(to_signed(957,16));
ROM(1263) <= std_logic_vector(to_signed(956,16));
ROM(1264) <= std_logic_vector(to_signed(955,16));
ROM(1265) <= std_logic_vector(to_signed(955,16));
ROM(1266) <= std_logic_vector(to_signed(954,16));
ROM(1267) <= std_logic_vector(to_signed(954,16));
ROM(1268) <= std_logic_vector(to_signed(953,16));
ROM(1269) <= std_logic_vector(to_signed(953,16));
ROM(1270) <= std_logic_vector(to_signed(952,16));
ROM(1271) <= std_logic_vector(to_signed(951,16));
ROM(1272) <= std_logic_vector(to_signed(951,16));
ROM(1273) <= std_logic_vector(to_signed(950,16));
ROM(1274) <= std_logic_vector(to_signed(950,16));
ROM(1275) <= std_logic_vector(to_signed(949,16));
ROM(1276) <= std_logic_vector(to_signed(948,16));
ROM(1277) <= std_logic_vector(to_signed(948,16));
ROM(1278) <= std_logic_vector(to_signed(947,16));
ROM(1279) <= std_logic_vector(to_signed(947,16));
ROM(1280) <= std_logic_vector(to_signed(946,16));
ROM(1281) <= std_logic_vector(to_signed(945,16));
ROM(1282) <= std_logic_vector(to_signed(945,16));
ROM(1283) <= std_logic_vector(to_signed(944,16));
ROM(1284) <= std_logic_vector(to_signed(944,16));
ROM(1285) <= std_logic_vector(to_signed(943,16));
ROM(1286) <= std_logic_vector(to_signed(942,16));
ROM(1287) <= std_logic_vector(to_signed(942,16));
ROM(1288) <= std_logic_vector(to_signed(941,16));
ROM(1289) <= std_logic_vector(to_signed(941,16));
ROM(1290) <= std_logic_vector(to_signed(940,16));
ROM(1291) <= std_logic_vector(to_signed(939,16));
ROM(1292) <= std_logic_vector(to_signed(939,16));
ROM(1293) <= std_logic_vector(to_signed(938,16));
ROM(1294) <= std_logic_vector(to_signed(937,16));
ROM(1295) <= std_logic_vector(to_signed(937,16));
ROM(1296) <= std_logic_vector(to_signed(936,16));
ROM(1297) <= std_logic_vector(to_signed(936,16));
ROM(1298) <= std_logic_vector(to_signed(935,16));
ROM(1299) <= std_logic_vector(to_signed(934,16));
ROM(1300) <= std_logic_vector(to_signed(934,16));
ROM(1301) <= std_logic_vector(to_signed(933,16));
ROM(1302) <= std_logic_vector(to_signed(932,16));
ROM(1303) <= std_logic_vector(to_signed(932,16));
ROM(1304) <= std_logic_vector(to_signed(931,16));
ROM(1305) <= std_logic_vector(to_signed(930,16));
ROM(1306) <= std_logic_vector(to_signed(930,16));
ROM(1307) <= std_logic_vector(to_signed(929,16));
ROM(1308) <= std_logic_vector(to_signed(928,16));
ROM(1309) <= std_logic_vector(to_signed(928,16));
ROM(1310) <= std_logic_vector(to_signed(927,16));
ROM(1311) <= std_logic_vector(to_signed(926,16));
ROM(1312) <= std_logic_vector(to_signed(926,16));
ROM(1313) <= std_logic_vector(to_signed(925,16));
ROM(1314) <= std_logic_vector(to_signed(924,16));
ROM(1315) <= std_logic_vector(to_signed(924,16));
ROM(1316) <= std_logic_vector(to_signed(923,16));
ROM(1317) <= std_logic_vector(to_signed(922,16));
ROM(1318) <= std_logic_vector(to_signed(922,16));
ROM(1319) <= std_logic_vector(to_signed(921,16));
ROM(1320) <= std_logic_vector(to_signed(920,16));
ROM(1321) <= std_logic_vector(to_signed(920,16));
ROM(1322) <= std_logic_vector(to_signed(919,16));
ROM(1323) <= std_logic_vector(to_signed(918,16));
ROM(1324) <= std_logic_vector(to_signed(917,16));
ROM(1325) <= std_logic_vector(to_signed(917,16));
ROM(1326) <= std_logic_vector(to_signed(916,16));
ROM(1327) <= std_logic_vector(to_signed(915,16));
ROM(1328) <= std_logic_vector(to_signed(915,16));
ROM(1329) <= std_logic_vector(to_signed(914,16));
ROM(1330) <= std_logic_vector(to_signed(913,16));
ROM(1331) <= std_logic_vector(to_signed(913,16));
ROM(1332) <= std_logic_vector(to_signed(912,16));
ROM(1333) <= std_logic_vector(to_signed(911,16));
ROM(1334) <= std_logic_vector(to_signed(910,16));
ROM(1335) <= std_logic_vector(to_signed(910,16));
ROM(1336) <= std_logic_vector(to_signed(909,16));
ROM(1337) <= std_logic_vector(to_signed(908,16));
ROM(1338) <= std_logic_vector(to_signed(907,16));
ROM(1339) <= std_logic_vector(to_signed(907,16));
ROM(1340) <= std_logic_vector(to_signed(906,16));
ROM(1341) <= std_logic_vector(to_signed(905,16));
ROM(1342) <= std_logic_vector(to_signed(905,16));
ROM(1343) <= std_logic_vector(to_signed(904,16));
ROM(1344) <= std_logic_vector(to_signed(903,16));
ROM(1345) <= std_logic_vector(to_signed(902,16));
ROM(1346) <= std_logic_vector(to_signed(902,16));
ROM(1347) <= std_logic_vector(to_signed(901,16));
ROM(1348) <= std_logic_vector(to_signed(900,16));
ROM(1349) <= std_logic_vector(to_signed(899,16));
ROM(1350) <= std_logic_vector(to_signed(899,16));
ROM(1351) <= std_logic_vector(to_signed(898,16));
ROM(1352) <= std_logic_vector(to_signed(897,16));
ROM(1353) <= std_logic_vector(to_signed(896,16));
ROM(1354) <= std_logic_vector(to_signed(896,16));
ROM(1355) <= std_logic_vector(to_signed(895,16));
ROM(1356) <= std_logic_vector(to_signed(894,16));
ROM(1357) <= std_logic_vector(to_signed(893,16));
ROM(1358) <= std_logic_vector(to_signed(893,16));
ROM(1359) <= std_logic_vector(to_signed(892,16));
ROM(1360) <= std_logic_vector(to_signed(891,16));
ROM(1361) <= std_logic_vector(to_signed(890,16));
ROM(1362) <= std_logic_vector(to_signed(889,16));
ROM(1363) <= std_logic_vector(to_signed(889,16));
ROM(1364) <= std_logic_vector(to_signed(888,16));
ROM(1365) <= std_logic_vector(to_signed(887,16));
ROM(1366) <= std_logic_vector(to_signed(886,16));
ROM(1367) <= std_logic_vector(to_signed(885,16));
ROM(1368) <= std_logic_vector(to_signed(885,16));
ROM(1369) <= std_logic_vector(to_signed(884,16));
ROM(1370) <= std_logic_vector(to_signed(883,16));
ROM(1371) <= std_logic_vector(to_signed(882,16));
ROM(1372) <= std_logic_vector(to_signed(882,16));
ROM(1373) <= std_logic_vector(to_signed(881,16));
ROM(1374) <= std_logic_vector(to_signed(880,16));
ROM(1375) <= std_logic_vector(to_signed(879,16));
ROM(1376) <= std_logic_vector(to_signed(878,16));
ROM(1377) <= std_logic_vector(to_signed(878,16));
ROM(1378) <= std_logic_vector(to_signed(877,16));
ROM(1379) <= std_logic_vector(to_signed(876,16));
ROM(1380) <= std_logic_vector(to_signed(875,16));
ROM(1381) <= std_logic_vector(to_signed(874,16));
ROM(1382) <= std_logic_vector(to_signed(873,16));
ROM(1383) <= std_logic_vector(to_signed(873,16));
ROM(1384) <= std_logic_vector(to_signed(872,16));
ROM(1385) <= std_logic_vector(to_signed(871,16));
ROM(1386) <= std_logic_vector(to_signed(870,16));
ROM(1387) <= std_logic_vector(to_signed(869,16));
ROM(1388) <= std_logic_vector(to_signed(868,16));
ROM(1389) <= std_logic_vector(to_signed(868,16));
ROM(1390) <= std_logic_vector(to_signed(867,16));
ROM(1391) <= std_logic_vector(to_signed(866,16));
ROM(1392) <= std_logic_vector(to_signed(865,16));
ROM(1393) <= std_logic_vector(to_signed(864,16));
ROM(1394) <= std_logic_vector(to_signed(863,16));
ROM(1395) <= std_logic_vector(to_signed(863,16));
ROM(1396) <= std_logic_vector(to_signed(862,16));
ROM(1397) <= std_logic_vector(to_signed(861,16));
ROM(1398) <= std_logic_vector(to_signed(860,16));
ROM(1399) <= std_logic_vector(to_signed(859,16));
ROM(1400) <= std_logic_vector(to_signed(858,16));
ROM(1401) <= std_logic_vector(to_signed(857,16));
ROM(1402) <= std_logic_vector(to_signed(857,16));
ROM(1403) <= std_logic_vector(to_signed(856,16));
ROM(1404) <= std_logic_vector(to_signed(855,16));
ROM(1405) <= std_logic_vector(to_signed(854,16));
ROM(1406) <= std_logic_vector(to_signed(853,16));
ROM(1407) <= std_logic_vector(to_signed(852,16));
ROM(1408) <= std_logic_vector(to_signed(851,16));
ROM(1409) <= std_logic_vector(to_signed(851,16));
ROM(1410) <= std_logic_vector(to_signed(850,16));
ROM(1411) <= std_logic_vector(to_signed(849,16));
ROM(1412) <= std_logic_vector(to_signed(848,16));
ROM(1413) <= std_logic_vector(to_signed(847,16));
ROM(1414) <= std_logic_vector(to_signed(846,16));
ROM(1415) <= std_logic_vector(to_signed(845,16));
ROM(1416) <= std_logic_vector(to_signed(844,16));
ROM(1417) <= std_logic_vector(to_signed(843,16));
ROM(1418) <= std_logic_vector(to_signed(843,16));
ROM(1419) <= std_logic_vector(to_signed(842,16));
ROM(1420) <= std_logic_vector(to_signed(841,16));
ROM(1421) <= std_logic_vector(to_signed(840,16));
ROM(1422) <= std_logic_vector(to_signed(839,16));
ROM(1423) <= std_logic_vector(to_signed(838,16));
ROM(1424) <= std_logic_vector(to_signed(837,16));
ROM(1425) <= std_logic_vector(to_signed(836,16));
ROM(1426) <= std_logic_vector(to_signed(835,16));
ROM(1427) <= std_logic_vector(to_signed(834,16));
ROM(1428) <= std_logic_vector(to_signed(834,16));
ROM(1429) <= std_logic_vector(to_signed(833,16));
ROM(1430) <= std_logic_vector(to_signed(832,16));
ROM(1431) <= std_logic_vector(to_signed(831,16));
ROM(1432) <= std_logic_vector(to_signed(830,16));
ROM(1433) <= std_logic_vector(to_signed(829,16));
ROM(1434) <= std_logic_vector(to_signed(828,16));
ROM(1435) <= std_logic_vector(to_signed(827,16));
ROM(1436) <= std_logic_vector(to_signed(826,16));
ROM(1437) <= std_logic_vector(to_signed(825,16));
ROM(1438) <= std_logic_vector(to_signed(824,16));
ROM(1439) <= std_logic_vector(to_signed(823,16));
ROM(1440) <= std_logic_vector(to_signed(822,16));
ROM(1441) <= std_logic_vector(to_signed(822,16));
ROM(1442) <= std_logic_vector(to_signed(821,16));
ROM(1443) <= std_logic_vector(to_signed(820,16));
ROM(1444) <= std_logic_vector(to_signed(819,16));
ROM(1445) <= std_logic_vector(to_signed(818,16));
ROM(1446) <= std_logic_vector(to_signed(817,16));
ROM(1447) <= std_logic_vector(to_signed(816,16));
ROM(1448) <= std_logic_vector(to_signed(815,16));
ROM(1449) <= std_logic_vector(to_signed(814,16));
ROM(1450) <= std_logic_vector(to_signed(813,16));
ROM(1451) <= std_logic_vector(to_signed(812,16));
ROM(1452) <= std_logic_vector(to_signed(811,16));
ROM(1453) <= std_logic_vector(to_signed(810,16));
ROM(1454) <= std_logic_vector(to_signed(809,16));
ROM(1455) <= std_logic_vector(to_signed(808,16));
ROM(1456) <= std_logic_vector(to_signed(807,16));
ROM(1457) <= std_logic_vector(to_signed(806,16));
ROM(1458) <= std_logic_vector(to_signed(805,16));
ROM(1459) <= std_logic_vector(to_signed(804,16));
ROM(1460) <= std_logic_vector(to_signed(803,16));
ROM(1461) <= std_logic_vector(to_signed(802,16));
ROM(1462) <= std_logic_vector(to_signed(801,16));
ROM(1463) <= std_logic_vector(to_signed(800,16));
ROM(1464) <= std_logic_vector(to_signed(799,16));
ROM(1465) <= std_logic_vector(to_signed(798,16));
ROM(1466) <= std_logic_vector(to_signed(798,16));
ROM(1467) <= std_logic_vector(to_signed(797,16));
ROM(1468) <= std_logic_vector(to_signed(796,16));
ROM(1469) <= std_logic_vector(to_signed(795,16));
ROM(1470) <= std_logic_vector(to_signed(794,16));
ROM(1471) <= std_logic_vector(to_signed(793,16));
ROM(1472) <= std_logic_vector(to_signed(792,16));
ROM(1473) <= std_logic_vector(to_signed(791,16));
ROM(1474) <= std_logic_vector(to_signed(790,16));
ROM(1475) <= std_logic_vector(to_signed(789,16));
ROM(1476) <= std_logic_vector(to_signed(788,16));
ROM(1477) <= std_logic_vector(to_signed(787,16));
ROM(1478) <= std_logic_vector(to_signed(786,16));
ROM(1479) <= std_logic_vector(to_signed(785,16));
ROM(1480) <= std_logic_vector(to_signed(784,16));
ROM(1481) <= std_logic_vector(to_signed(783,16));
ROM(1482) <= std_logic_vector(to_signed(782,16));
ROM(1483) <= std_logic_vector(to_signed(780,16));
ROM(1484) <= std_logic_vector(to_signed(779,16));
ROM(1485) <= std_logic_vector(to_signed(778,16));
ROM(1486) <= std_logic_vector(to_signed(777,16));
ROM(1487) <= std_logic_vector(to_signed(776,16));
ROM(1488) <= std_logic_vector(to_signed(775,16));
ROM(1489) <= std_logic_vector(to_signed(774,16));
ROM(1490) <= std_logic_vector(to_signed(773,16));
ROM(1491) <= std_logic_vector(to_signed(772,16));
ROM(1492) <= std_logic_vector(to_signed(771,16));
ROM(1493) <= std_logic_vector(to_signed(770,16));
ROM(1494) <= std_logic_vector(to_signed(769,16));
ROM(1495) <= std_logic_vector(to_signed(768,16));
ROM(1496) <= std_logic_vector(to_signed(767,16));
ROM(1497) <= std_logic_vector(to_signed(766,16));
ROM(1498) <= std_logic_vector(to_signed(765,16));
ROM(1499) <= std_logic_vector(to_signed(764,16));
ROM(1500) <= std_logic_vector(to_signed(763,16));
ROM(1501) <= std_logic_vector(to_signed(762,16));
ROM(1502) <= std_logic_vector(to_signed(761,16));
ROM(1503) <= std_logic_vector(to_signed(760,16));
ROM(1504) <= std_logic_vector(to_signed(759,16));
ROM(1505) <= std_logic_vector(to_signed(758,16));
ROM(1506) <= std_logic_vector(to_signed(757,16));
ROM(1507) <= std_logic_vector(to_signed(756,16));
ROM(1508) <= std_logic_vector(to_signed(755,16));
ROM(1509) <= std_logic_vector(to_signed(753,16));
ROM(1510) <= std_logic_vector(to_signed(752,16));
ROM(1511) <= std_logic_vector(to_signed(751,16));
ROM(1512) <= std_logic_vector(to_signed(750,16));
ROM(1513) <= std_logic_vector(to_signed(749,16));
ROM(1514) <= std_logic_vector(to_signed(748,16));
ROM(1515) <= std_logic_vector(to_signed(747,16));
ROM(1516) <= std_logic_vector(to_signed(746,16));
ROM(1517) <= std_logic_vector(to_signed(745,16));
ROM(1518) <= std_logic_vector(to_signed(744,16));
ROM(1519) <= std_logic_vector(to_signed(743,16));
ROM(1520) <= std_logic_vector(to_signed(742,16));
ROM(1521) <= std_logic_vector(to_signed(741,16));
ROM(1522) <= std_logic_vector(to_signed(739,16));
ROM(1523) <= std_logic_vector(to_signed(738,16));
ROM(1524) <= std_logic_vector(to_signed(737,16));
ROM(1525) <= std_logic_vector(to_signed(736,16));
ROM(1526) <= std_logic_vector(to_signed(735,16));
ROM(1527) <= std_logic_vector(to_signed(734,16));
ROM(1528) <= std_logic_vector(to_signed(733,16));
ROM(1529) <= std_logic_vector(to_signed(732,16));
ROM(1530) <= std_logic_vector(to_signed(731,16));
ROM(1531) <= std_logic_vector(to_signed(730,16));
ROM(1532) <= std_logic_vector(to_signed(729,16));
ROM(1533) <= std_logic_vector(to_signed(727,16));
ROM(1534) <= std_logic_vector(to_signed(726,16));
ROM(1535) <= std_logic_vector(to_signed(725,16));
ROM(1536) <= std_logic_vector(to_signed(724,16));
ROM(1537) <= std_logic_vector(to_signed(723,16));
ROM(1538) <= std_logic_vector(to_signed(722,16));
ROM(1539) <= std_logic_vector(to_signed(721,16));
ROM(1540) <= std_logic_vector(to_signed(720,16));
ROM(1541) <= std_logic_vector(to_signed(719,16));
ROM(1542) <= std_logic_vector(to_signed(717,16));
ROM(1543) <= std_logic_vector(to_signed(716,16));
ROM(1544) <= std_logic_vector(to_signed(715,16));
ROM(1545) <= std_logic_vector(to_signed(714,16));
ROM(1546) <= std_logic_vector(to_signed(713,16));
ROM(1547) <= std_logic_vector(to_signed(712,16));
ROM(1548) <= std_logic_vector(to_signed(711,16));
ROM(1549) <= std_logic_vector(to_signed(709,16));
ROM(1550) <= std_logic_vector(to_signed(708,16));
ROM(1551) <= std_logic_vector(to_signed(707,16));
ROM(1552) <= std_logic_vector(to_signed(706,16));
ROM(1553) <= std_logic_vector(to_signed(705,16));
ROM(1554) <= std_logic_vector(to_signed(704,16));
ROM(1555) <= std_logic_vector(to_signed(703,16));
ROM(1556) <= std_logic_vector(to_signed(702,16));
ROM(1557) <= std_logic_vector(to_signed(700,16));
ROM(1558) <= std_logic_vector(to_signed(699,16));
ROM(1559) <= std_logic_vector(to_signed(698,16));
ROM(1560) <= std_logic_vector(to_signed(697,16));
ROM(1561) <= std_logic_vector(to_signed(696,16));
ROM(1562) <= std_logic_vector(to_signed(695,16));
ROM(1563) <= std_logic_vector(to_signed(693,16));
ROM(1564) <= std_logic_vector(to_signed(692,16));
ROM(1565) <= std_logic_vector(to_signed(691,16));
ROM(1566) <= std_logic_vector(to_signed(690,16));
ROM(1567) <= std_logic_vector(to_signed(689,16));
ROM(1568) <= std_logic_vector(to_signed(688,16));
ROM(1569) <= std_logic_vector(to_signed(687,16));
ROM(1570) <= std_logic_vector(to_signed(685,16));
ROM(1571) <= std_logic_vector(to_signed(684,16));
ROM(1572) <= std_logic_vector(to_signed(683,16));
ROM(1573) <= std_logic_vector(to_signed(682,16));
ROM(1574) <= std_logic_vector(to_signed(681,16));
ROM(1575) <= std_logic_vector(to_signed(679,16));
ROM(1576) <= std_logic_vector(to_signed(678,16));
ROM(1577) <= std_logic_vector(to_signed(677,16));
ROM(1578) <= std_logic_vector(to_signed(676,16));
ROM(1579) <= std_logic_vector(to_signed(675,16));
ROM(1580) <= std_logic_vector(to_signed(674,16));
ROM(1581) <= std_logic_vector(to_signed(672,16));
ROM(1582) <= std_logic_vector(to_signed(671,16));
ROM(1583) <= std_logic_vector(to_signed(670,16));
ROM(1584) <= std_logic_vector(to_signed(669,16));
ROM(1585) <= std_logic_vector(to_signed(668,16));
ROM(1586) <= std_logic_vector(to_signed(666,16));
ROM(1587) <= std_logic_vector(to_signed(665,16));
ROM(1588) <= std_logic_vector(to_signed(664,16));
ROM(1589) <= std_logic_vector(to_signed(663,16));
ROM(1590) <= std_logic_vector(to_signed(662,16));
ROM(1591) <= std_logic_vector(to_signed(660,16));
ROM(1592) <= std_logic_vector(to_signed(659,16));
ROM(1593) <= std_logic_vector(to_signed(658,16));
ROM(1594) <= std_logic_vector(to_signed(657,16));
ROM(1595) <= std_logic_vector(to_signed(656,16));
ROM(1596) <= std_logic_vector(to_signed(654,16));
ROM(1597) <= std_logic_vector(to_signed(653,16));
ROM(1598) <= std_logic_vector(to_signed(652,16));
ROM(1599) <= std_logic_vector(to_signed(651,16));
ROM(1600) <= std_logic_vector(to_signed(650,16));
ROM(1601) <= std_logic_vector(to_signed(648,16));
ROM(1602) <= std_logic_vector(to_signed(647,16));
ROM(1603) <= std_logic_vector(to_signed(646,16));
ROM(1604) <= std_logic_vector(to_signed(645,16));
ROM(1605) <= std_logic_vector(to_signed(644,16));
ROM(1606) <= std_logic_vector(to_signed(642,16));
ROM(1607) <= std_logic_vector(to_signed(641,16));
ROM(1608) <= std_logic_vector(to_signed(640,16));
ROM(1609) <= std_logic_vector(to_signed(639,16));
ROM(1610) <= std_logic_vector(to_signed(637,16));
ROM(1611) <= std_logic_vector(to_signed(636,16));
ROM(1612) <= std_logic_vector(to_signed(635,16));
ROM(1613) <= std_logic_vector(to_signed(634,16));
ROM(1614) <= std_logic_vector(to_signed(632,16));
ROM(1615) <= std_logic_vector(to_signed(631,16));
ROM(1616) <= std_logic_vector(to_signed(630,16));
ROM(1617) <= std_logic_vector(to_signed(629,16));
ROM(1618) <= std_logic_vector(to_signed(628,16));
ROM(1619) <= std_logic_vector(to_signed(626,16));
ROM(1620) <= std_logic_vector(to_signed(625,16));
ROM(1621) <= std_logic_vector(to_signed(624,16));
ROM(1622) <= std_logic_vector(to_signed(623,16));
ROM(1623) <= std_logic_vector(to_signed(621,16));
ROM(1624) <= std_logic_vector(to_signed(620,16));
ROM(1625) <= std_logic_vector(to_signed(619,16));
ROM(1626) <= std_logic_vector(to_signed(618,16));
ROM(1627) <= std_logic_vector(to_signed(616,16));
ROM(1628) <= std_logic_vector(to_signed(615,16));
ROM(1629) <= std_logic_vector(to_signed(614,16));
ROM(1630) <= std_logic_vector(to_signed(613,16));
ROM(1631) <= std_logic_vector(to_signed(611,16));
ROM(1632) <= std_logic_vector(to_signed(610,16));
ROM(1633) <= std_logic_vector(to_signed(609,16));
ROM(1634) <= std_logic_vector(to_signed(607,16));
ROM(1635) <= std_logic_vector(to_signed(606,16));
ROM(1636) <= std_logic_vector(to_signed(605,16));
ROM(1637) <= std_logic_vector(to_signed(604,16));
ROM(1638) <= std_logic_vector(to_signed(602,16));
ROM(1639) <= std_logic_vector(to_signed(601,16));
ROM(1640) <= std_logic_vector(to_signed(600,16));
ROM(1641) <= std_logic_vector(to_signed(599,16));
ROM(1642) <= std_logic_vector(to_signed(597,16));
ROM(1643) <= std_logic_vector(to_signed(596,16));
ROM(1644) <= std_logic_vector(to_signed(595,16));
ROM(1645) <= std_logic_vector(to_signed(593,16));
ROM(1646) <= std_logic_vector(to_signed(592,16));
ROM(1647) <= std_logic_vector(to_signed(591,16));
ROM(1648) <= std_logic_vector(to_signed(590,16));
ROM(1649) <= std_logic_vector(to_signed(588,16));
ROM(1650) <= std_logic_vector(to_signed(587,16));
ROM(1651) <= std_logic_vector(to_signed(586,16));
ROM(1652) <= std_logic_vector(to_signed(584,16));
ROM(1653) <= std_logic_vector(to_signed(583,16));
ROM(1654) <= std_logic_vector(to_signed(582,16));
ROM(1655) <= std_logic_vector(to_signed(581,16));
ROM(1656) <= std_logic_vector(to_signed(579,16));
ROM(1657) <= std_logic_vector(to_signed(578,16));
ROM(1658) <= std_logic_vector(to_signed(577,16));
ROM(1659) <= std_logic_vector(to_signed(575,16));
ROM(1660) <= std_logic_vector(to_signed(574,16));
ROM(1661) <= std_logic_vector(to_signed(573,16));
ROM(1662) <= std_logic_vector(to_signed(572,16));
ROM(1663) <= std_logic_vector(to_signed(570,16));
ROM(1664) <= std_logic_vector(to_signed(569,16));
ROM(1665) <= std_logic_vector(to_signed(568,16));
ROM(1666) <= std_logic_vector(to_signed(566,16));
ROM(1667) <= std_logic_vector(to_signed(565,16));
ROM(1668) <= std_logic_vector(to_signed(564,16));
ROM(1669) <= std_logic_vector(to_signed(562,16));
ROM(1670) <= std_logic_vector(to_signed(561,16));
ROM(1671) <= std_logic_vector(to_signed(560,16));
ROM(1672) <= std_logic_vector(to_signed(558,16));
ROM(1673) <= std_logic_vector(to_signed(557,16));
ROM(1674) <= std_logic_vector(to_signed(556,16));
ROM(1675) <= std_logic_vector(to_signed(554,16));
ROM(1676) <= std_logic_vector(to_signed(553,16));
ROM(1677) <= std_logic_vector(to_signed(552,16));
ROM(1678) <= std_logic_vector(to_signed(550,16));
ROM(1679) <= std_logic_vector(to_signed(549,16));
ROM(1680) <= std_logic_vector(to_signed(548,16));
ROM(1681) <= std_logic_vector(to_signed(547,16));
ROM(1682) <= std_logic_vector(to_signed(545,16));
ROM(1683) <= std_logic_vector(to_signed(544,16));
ROM(1684) <= std_logic_vector(to_signed(543,16));
ROM(1685) <= std_logic_vector(to_signed(541,16));
ROM(1686) <= std_logic_vector(to_signed(540,16));
ROM(1687) <= std_logic_vector(to_signed(539,16));
ROM(1688) <= std_logic_vector(to_signed(537,16));
ROM(1689) <= std_logic_vector(to_signed(536,16));
ROM(1690) <= std_logic_vector(to_signed(535,16));
ROM(1691) <= std_logic_vector(to_signed(533,16));
ROM(1692) <= std_logic_vector(to_signed(532,16));
ROM(1693) <= std_logic_vector(to_signed(530,16));
ROM(1694) <= std_logic_vector(to_signed(529,16));
ROM(1695) <= std_logic_vector(to_signed(528,16));
ROM(1696) <= std_logic_vector(to_signed(526,16));
ROM(1697) <= std_logic_vector(to_signed(525,16));
ROM(1698) <= std_logic_vector(to_signed(524,16));
ROM(1699) <= std_logic_vector(to_signed(522,16));
ROM(1700) <= std_logic_vector(to_signed(521,16));
ROM(1701) <= std_logic_vector(to_signed(520,16));
ROM(1702) <= std_logic_vector(to_signed(518,16));
ROM(1703) <= std_logic_vector(to_signed(517,16));
ROM(1704) <= std_logic_vector(to_signed(516,16));
ROM(1705) <= std_logic_vector(to_signed(514,16));
ROM(1706) <= std_logic_vector(to_signed(513,16));
ROM(1707) <= std_logic_vector(to_signed(512,16));
ROM(1708) <= std_logic_vector(to_signed(510,16));
ROM(1709) <= std_logic_vector(to_signed(509,16));
ROM(1710) <= std_logic_vector(to_signed(507,16));
ROM(1711) <= std_logic_vector(to_signed(506,16));
ROM(1712) <= std_logic_vector(to_signed(505,16));
ROM(1713) <= std_logic_vector(to_signed(503,16));
ROM(1714) <= std_logic_vector(to_signed(502,16));
ROM(1715) <= std_logic_vector(to_signed(501,16));
ROM(1716) <= std_logic_vector(to_signed(499,16));
ROM(1717) <= std_logic_vector(to_signed(498,16));
ROM(1718) <= std_logic_vector(to_signed(497,16));
ROM(1719) <= std_logic_vector(to_signed(495,16));
ROM(1720) <= std_logic_vector(to_signed(494,16));
ROM(1721) <= std_logic_vector(to_signed(492,16));
ROM(1722) <= std_logic_vector(to_signed(491,16));
ROM(1723) <= std_logic_vector(to_signed(490,16));
ROM(1724) <= std_logic_vector(to_signed(488,16));
ROM(1725) <= std_logic_vector(to_signed(487,16));
ROM(1726) <= std_logic_vector(to_signed(485,16));
ROM(1727) <= std_logic_vector(to_signed(484,16));
ROM(1728) <= std_logic_vector(to_signed(483,16));
ROM(1729) <= std_logic_vector(to_signed(481,16));
ROM(1730) <= std_logic_vector(to_signed(480,16));
ROM(1731) <= std_logic_vector(to_signed(479,16));
ROM(1732) <= std_logic_vector(to_signed(477,16));
ROM(1733) <= std_logic_vector(to_signed(476,16));
ROM(1734) <= std_logic_vector(to_signed(474,16));
ROM(1735) <= std_logic_vector(to_signed(473,16));
ROM(1736) <= std_logic_vector(to_signed(472,16));
ROM(1737) <= std_logic_vector(to_signed(470,16));
ROM(1738) <= std_logic_vector(to_signed(469,16));
ROM(1739) <= std_logic_vector(to_signed(467,16));
ROM(1740) <= std_logic_vector(to_signed(466,16));
ROM(1741) <= std_logic_vector(to_signed(465,16));
ROM(1742) <= std_logic_vector(to_signed(463,16));
ROM(1743) <= std_logic_vector(to_signed(462,16));
ROM(1744) <= std_logic_vector(to_signed(460,16));
ROM(1745) <= std_logic_vector(to_signed(459,16));
ROM(1746) <= std_logic_vector(to_signed(458,16));
ROM(1747) <= std_logic_vector(to_signed(456,16));
ROM(1748) <= std_logic_vector(to_signed(455,16));
ROM(1749) <= std_logic_vector(to_signed(453,16));
ROM(1750) <= std_logic_vector(to_signed(452,16));
ROM(1751) <= std_logic_vector(to_signed(451,16));
ROM(1752) <= std_logic_vector(to_signed(449,16));
ROM(1753) <= std_logic_vector(to_signed(448,16));
ROM(1754) <= std_logic_vector(to_signed(446,16));
ROM(1755) <= std_logic_vector(to_signed(445,16));
ROM(1756) <= std_logic_vector(to_signed(443,16));
ROM(1757) <= std_logic_vector(to_signed(442,16));
ROM(1758) <= std_logic_vector(to_signed(441,16));
ROM(1759) <= std_logic_vector(to_signed(439,16));
ROM(1760) <= std_logic_vector(to_signed(438,16));
ROM(1761) <= std_logic_vector(to_signed(436,16));
ROM(1762) <= std_logic_vector(to_signed(435,16));
ROM(1763) <= std_logic_vector(to_signed(434,16));
ROM(1764) <= std_logic_vector(to_signed(432,16));
ROM(1765) <= std_logic_vector(to_signed(431,16));
ROM(1766) <= std_logic_vector(to_signed(429,16));
ROM(1767) <= std_logic_vector(to_signed(428,16));
ROM(1768) <= std_logic_vector(to_signed(426,16));
ROM(1769) <= std_logic_vector(to_signed(425,16));
ROM(1770) <= std_logic_vector(to_signed(424,16));
ROM(1771) <= std_logic_vector(to_signed(422,16));
ROM(1772) <= std_logic_vector(to_signed(421,16));
ROM(1773) <= std_logic_vector(to_signed(419,16));
ROM(1774) <= std_logic_vector(to_signed(418,16));
ROM(1775) <= std_logic_vector(to_signed(416,16));
ROM(1776) <= std_logic_vector(to_signed(415,16));
ROM(1777) <= std_logic_vector(to_signed(414,16));
ROM(1778) <= std_logic_vector(to_signed(412,16));
ROM(1779) <= std_logic_vector(to_signed(411,16));
ROM(1780) <= std_logic_vector(to_signed(409,16));
ROM(1781) <= std_logic_vector(to_signed(408,16));
ROM(1782) <= std_logic_vector(to_signed(406,16));
ROM(1783) <= std_logic_vector(to_signed(405,16));
ROM(1784) <= std_logic_vector(to_signed(403,16));
ROM(1785) <= std_logic_vector(to_signed(402,16));
ROM(1786) <= std_logic_vector(to_signed(401,16));
ROM(1787) <= std_logic_vector(to_signed(399,16));
ROM(1788) <= std_logic_vector(to_signed(398,16));
ROM(1789) <= std_logic_vector(to_signed(396,16));
ROM(1790) <= std_logic_vector(to_signed(395,16));
ROM(1791) <= std_logic_vector(to_signed(393,16));
ROM(1792) <= std_logic_vector(to_signed(392,16));
ROM(1793) <= std_logic_vector(to_signed(390,16));
ROM(1794) <= std_logic_vector(to_signed(389,16));
ROM(1795) <= std_logic_vector(to_signed(388,16));
ROM(1796) <= std_logic_vector(to_signed(386,16));
ROM(1797) <= std_logic_vector(to_signed(385,16));
ROM(1798) <= std_logic_vector(to_signed(383,16));
ROM(1799) <= std_logic_vector(to_signed(382,16));
ROM(1800) <= std_logic_vector(to_signed(380,16));
ROM(1801) <= std_logic_vector(to_signed(379,16));
ROM(1802) <= std_logic_vector(to_signed(377,16));
ROM(1803) <= std_logic_vector(to_signed(376,16));
ROM(1804) <= std_logic_vector(to_signed(374,16));
ROM(1805) <= std_logic_vector(to_signed(373,16));
ROM(1806) <= std_logic_vector(to_signed(371,16));
ROM(1807) <= std_logic_vector(to_signed(370,16));
ROM(1808) <= std_logic_vector(to_signed(369,16));
ROM(1809) <= std_logic_vector(to_signed(367,16));
ROM(1810) <= std_logic_vector(to_signed(366,16));
ROM(1811) <= std_logic_vector(to_signed(364,16));
ROM(1812) <= std_logic_vector(to_signed(363,16));
ROM(1813) <= std_logic_vector(to_signed(361,16));
ROM(1814) <= std_logic_vector(to_signed(360,16));
ROM(1815) <= std_logic_vector(to_signed(358,16));
ROM(1816) <= std_logic_vector(to_signed(357,16));
ROM(1817) <= std_logic_vector(to_signed(355,16));
ROM(1818) <= std_logic_vector(to_signed(354,16));
ROM(1819) <= std_logic_vector(to_signed(352,16));
ROM(1820) <= std_logic_vector(to_signed(351,16));
ROM(1821) <= std_logic_vector(to_signed(349,16));
ROM(1822) <= std_logic_vector(to_signed(348,16));
ROM(1823) <= std_logic_vector(to_signed(346,16));
ROM(1824) <= std_logic_vector(to_signed(345,16));
ROM(1825) <= std_logic_vector(to_signed(343,16));
ROM(1826) <= std_logic_vector(to_signed(342,16));
ROM(1827) <= std_logic_vector(to_signed(341,16));
ROM(1828) <= std_logic_vector(to_signed(339,16));
ROM(1829) <= std_logic_vector(to_signed(338,16));
ROM(1830) <= std_logic_vector(to_signed(336,16));
ROM(1831) <= std_logic_vector(to_signed(335,16));
ROM(1832) <= std_logic_vector(to_signed(333,16));
ROM(1833) <= std_logic_vector(to_signed(332,16));
ROM(1834) <= std_logic_vector(to_signed(330,16));
ROM(1835) <= std_logic_vector(to_signed(329,16));
ROM(1836) <= std_logic_vector(to_signed(327,16));
ROM(1837) <= std_logic_vector(to_signed(326,16));
ROM(1838) <= std_logic_vector(to_signed(324,16));
ROM(1839) <= std_logic_vector(to_signed(323,16));
ROM(1840) <= std_logic_vector(to_signed(321,16));
ROM(1841) <= std_logic_vector(to_signed(320,16));
ROM(1842) <= std_logic_vector(to_signed(318,16));
ROM(1843) <= std_logic_vector(to_signed(317,16));
ROM(1844) <= std_logic_vector(to_signed(315,16));
ROM(1845) <= std_logic_vector(to_signed(314,16));
ROM(1846) <= std_logic_vector(to_signed(312,16));
ROM(1847) <= std_logic_vector(to_signed(311,16));
ROM(1848) <= std_logic_vector(to_signed(309,16));
ROM(1849) <= std_logic_vector(to_signed(308,16));
ROM(1850) <= std_logic_vector(to_signed(306,16));
ROM(1851) <= std_logic_vector(to_signed(305,16));
ROM(1852) <= std_logic_vector(to_signed(303,16));
ROM(1853) <= std_logic_vector(to_signed(302,16));
ROM(1854) <= std_logic_vector(to_signed(300,16));
ROM(1855) <= std_logic_vector(to_signed(299,16));
ROM(1856) <= std_logic_vector(to_signed(297,16));
ROM(1857) <= std_logic_vector(to_signed(296,16));
ROM(1858) <= std_logic_vector(to_signed(294,16));
ROM(1859) <= std_logic_vector(to_signed(293,16));
ROM(1860) <= std_logic_vector(to_signed(291,16));
ROM(1861) <= std_logic_vector(to_signed(290,16));
ROM(1862) <= std_logic_vector(to_signed(288,16));
ROM(1863) <= std_logic_vector(to_signed(287,16));
ROM(1864) <= std_logic_vector(to_signed(285,16));
ROM(1865) <= std_logic_vector(to_signed(284,16));
ROM(1866) <= std_logic_vector(to_signed(282,16));
ROM(1867) <= std_logic_vector(to_signed(281,16));
ROM(1868) <= std_logic_vector(to_signed(279,16));
ROM(1869) <= std_logic_vector(to_signed(278,16));
ROM(1870) <= std_logic_vector(to_signed(276,16));
ROM(1871) <= std_logic_vector(to_signed(275,16));
ROM(1872) <= std_logic_vector(to_signed(273,16));
ROM(1873) <= std_logic_vector(to_signed(272,16));
ROM(1874) <= std_logic_vector(to_signed(270,16));
ROM(1875) <= std_logic_vector(to_signed(269,16));
ROM(1876) <= std_logic_vector(to_signed(267,16));
ROM(1877) <= std_logic_vector(to_signed(266,16));
ROM(1878) <= std_logic_vector(to_signed(264,16));
ROM(1879) <= std_logic_vector(to_signed(263,16));
ROM(1880) <= std_logic_vector(to_signed(261,16));
ROM(1881) <= std_logic_vector(to_signed(259,16));
ROM(1882) <= std_logic_vector(to_signed(258,16));
ROM(1883) <= std_logic_vector(to_signed(256,16));
ROM(1884) <= std_logic_vector(to_signed(255,16));
ROM(1885) <= std_logic_vector(to_signed(253,16));
ROM(1886) <= std_logic_vector(to_signed(252,16));
ROM(1887) <= std_logic_vector(to_signed(250,16));
ROM(1888) <= std_logic_vector(to_signed(249,16));
ROM(1889) <= std_logic_vector(to_signed(247,16));
ROM(1890) <= std_logic_vector(to_signed(246,16));
ROM(1891) <= std_logic_vector(to_signed(244,16));
ROM(1892) <= std_logic_vector(to_signed(243,16));
ROM(1893) <= std_logic_vector(to_signed(241,16));
ROM(1894) <= std_logic_vector(to_signed(240,16));
ROM(1895) <= std_logic_vector(to_signed(238,16));
ROM(1896) <= std_logic_vector(to_signed(237,16));
ROM(1897) <= std_logic_vector(to_signed(235,16));
ROM(1898) <= std_logic_vector(to_signed(234,16));
ROM(1899) <= std_logic_vector(to_signed(232,16));
ROM(1900) <= std_logic_vector(to_signed(230,16));
ROM(1901) <= std_logic_vector(to_signed(229,16));
ROM(1902) <= std_logic_vector(to_signed(227,16));
ROM(1903) <= std_logic_vector(to_signed(226,16));
ROM(1904) <= std_logic_vector(to_signed(224,16));
ROM(1905) <= std_logic_vector(to_signed(223,16));
ROM(1906) <= std_logic_vector(to_signed(221,16));
ROM(1907) <= std_logic_vector(to_signed(220,16));
ROM(1908) <= std_logic_vector(to_signed(218,16));
ROM(1909) <= std_logic_vector(to_signed(217,16));
ROM(1910) <= std_logic_vector(to_signed(215,16));
ROM(1911) <= std_logic_vector(to_signed(214,16));
ROM(1912) <= std_logic_vector(to_signed(212,16));
ROM(1913) <= std_logic_vector(to_signed(211,16));
ROM(1914) <= std_logic_vector(to_signed(209,16));
ROM(1915) <= std_logic_vector(to_signed(207,16));
ROM(1916) <= std_logic_vector(to_signed(206,16));
ROM(1917) <= std_logic_vector(to_signed(204,16));
ROM(1918) <= std_logic_vector(to_signed(203,16));
ROM(1919) <= std_logic_vector(to_signed(201,16));
ROM(1920) <= std_logic_vector(to_signed(200,16));
ROM(1921) <= std_logic_vector(to_signed(198,16));
ROM(1922) <= std_logic_vector(to_signed(197,16));
ROM(1923) <= std_logic_vector(to_signed(195,16));
ROM(1924) <= std_logic_vector(to_signed(194,16));
ROM(1925) <= std_logic_vector(to_signed(192,16));
ROM(1926) <= std_logic_vector(to_signed(191,16));
ROM(1927) <= std_logic_vector(to_signed(189,16));
ROM(1928) <= std_logic_vector(to_signed(187,16));
ROM(1929) <= std_logic_vector(to_signed(186,16));
ROM(1930) <= std_logic_vector(to_signed(184,16));
ROM(1931) <= std_logic_vector(to_signed(183,16));
ROM(1932) <= std_logic_vector(to_signed(181,16));
ROM(1933) <= std_logic_vector(to_signed(180,16));
ROM(1934) <= std_logic_vector(to_signed(178,16));
ROM(1935) <= std_logic_vector(to_signed(177,16));
ROM(1936) <= std_logic_vector(to_signed(175,16));
ROM(1937) <= std_logic_vector(to_signed(174,16));
ROM(1938) <= std_logic_vector(to_signed(172,16));
ROM(1939) <= std_logic_vector(to_signed(170,16));
ROM(1940) <= std_logic_vector(to_signed(169,16));
ROM(1941) <= std_logic_vector(to_signed(167,16));
ROM(1942) <= std_logic_vector(to_signed(166,16));
ROM(1943) <= std_logic_vector(to_signed(164,16));
ROM(1944) <= std_logic_vector(to_signed(163,16));
ROM(1945) <= std_logic_vector(to_signed(161,16));
ROM(1946) <= std_logic_vector(to_signed(160,16));
ROM(1947) <= std_logic_vector(to_signed(158,16));
ROM(1948) <= std_logic_vector(to_signed(156,16));
ROM(1949) <= std_logic_vector(to_signed(155,16));
ROM(1950) <= std_logic_vector(to_signed(153,16));
ROM(1951) <= std_logic_vector(to_signed(152,16));
ROM(1952) <= std_logic_vector(to_signed(150,16));
ROM(1953) <= std_logic_vector(to_signed(149,16));
ROM(1954) <= std_logic_vector(to_signed(147,16));
ROM(1955) <= std_logic_vector(to_signed(146,16));
ROM(1956) <= std_logic_vector(to_signed(144,16));
ROM(1957) <= std_logic_vector(to_signed(142,16));
ROM(1958) <= std_logic_vector(to_signed(141,16));
ROM(1959) <= std_logic_vector(to_signed(139,16));
ROM(1960) <= std_logic_vector(to_signed(138,16));
ROM(1961) <= std_logic_vector(to_signed(136,16));
ROM(1962) <= std_logic_vector(to_signed(135,16));
ROM(1963) <= std_logic_vector(to_signed(133,16));
ROM(1964) <= std_logic_vector(to_signed(132,16));
ROM(1965) <= std_logic_vector(to_signed(130,16));
ROM(1966) <= std_logic_vector(to_signed(128,16));
ROM(1967) <= std_logic_vector(to_signed(127,16));
ROM(1968) <= std_logic_vector(to_signed(125,16));
ROM(1969) <= std_logic_vector(to_signed(124,16));
ROM(1970) <= std_logic_vector(to_signed(122,16));
ROM(1971) <= std_logic_vector(to_signed(121,16));
ROM(1972) <= std_logic_vector(to_signed(119,16));
ROM(1973) <= std_logic_vector(to_signed(118,16));
ROM(1974) <= std_logic_vector(to_signed(116,16));
ROM(1975) <= std_logic_vector(to_signed(114,16));
ROM(1976) <= std_logic_vector(to_signed(113,16));
ROM(1977) <= std_logic_vector(to_signed(111,16));
ROM(1978) <= std_logic_vector(to_signed(110,16));
ROM(1979) <= std_logic_vector(to_signed(108,16));
ROM(1980) <= std_logic_vector(to_signed(107,16));
ROM(1981) <= std_logic_vector(to_signed(105,16));
ROM(1982) <= std_logic_vector(to_signed(103,16));
ROM(1983) <= std_logic_vector(to_signed(102,16));
ROM(1984) <= std_logic_vector(to_signed(100,16));
ROM(1985) <= std_logic_vector(to_signed(99,16));
ROM(1986) <= std_logic_vector(to_signed(97,16));
ROM(1987) <= std_logic_vector(to_signed(96,16));
ROM(1988) <= std_logic_vector(to_signed(94,16));
ROM(1989) <= std_logic_vector(to_signed(93,16));
ROM(1990) <= std_logic_vector(to_signed(91,16));
ROM(1991) <= std_logic_vector(to_signed(89,16));
ROM(1992) <= std_logic_vector(to_signed(88,16));
ROM(1993) <= std_logic_vector(to_signed(86,16));
ROM(1994) <= std_logic_vector(to_signed(85,16));
ROM(1995) <= std_logic_vector(to_signed(83,16));
ROM(1996) <= std_logic_vector(to_signed(82,16));
ROM(1997) <= std_logic_vector(to_signed(80,16));
ROM(1998) <= std_logic_vector(to_signed(78,16));
ROM(1999) <= std_logic_vector(to_signed(77,16));
ROM(2000) <= std_logic_vector(to_signed(75,16));
ROM(2001) <= std_logic_vector(to_signed(74,16));
ROM(2002) <= std_logic_vector(to_signed(72,16));
ROM(2003) <= std_logic_vector(to_signed(71,16));
ROM(2004) <= std_logic_vector(to_signed(69,16));
ROM(2005) <= std_logic_vector(to_signed(67,16));
ROM(2006) <= std_logic_vector(to_signed(66,16));
ROM(2007) <= std_logic_vector(to_signed(64,16));
ROM(2008) <= std_logic_vector(to_signed(63,16));
ROM(2009) <= std_logic_vector(to_signed(61,16));
ROM(2010) <= std_logic_vector(to_signed(60,16));
ROM(2011) <= std_logic_vector(to_signed(58,16));
ROM(2012) <= std_logic_vector(to_signed(57,16));
ROM(2013) <= std_logic_vector(to_signed(55,16));
ROM(2014) <= std_logic_vector(to_signed(53,16));
ROM(2015) <= std_logic_vector(to_signed(52,16));
ROM(2016) <= std_logic_vector(to_signed(50,16));
ROM(2017) <= std_logic_vector(to_signed(49,16));
ROM(2018) <= std_logic_vector(to_signed(47,16));
ROM(2019) <= std_logic_vector(to_signed(46,16));
ROM(2020) <= std_logic_vector(to_signed(44,16));
ROM(2021) <= std_logic_vector(to_signed(42,16));
ROM(2022) <= std_logic_vector(to_signed(41,16));
ROM(2023) <= std_logic_vector(to_signed(39,16));
ROM(2024) <= std_logic_vector(to_signed(38,16));
ROM(2025) <= std_logic_vector(to_signed(36,16));
ROM(2026) <= std_logic_vector(to_signed(35,16));
ROM(2027) <= std_logic_vector(to_signed(33,16));
ROM(2028) <= std_logic_vector(to_signed(31,16));
ROM(2029) <= std_logic_vector(to_signed(30,16));
ROM(2030) <= std_logic_vector(to_signed(28,16));
ROM(2031) <= std_logic_vector(to_signed(27,16));
ROM(2032) <= std_logic_vector(to_signed(25,16));
ROM(2033) <= std_logic_vector(to_signed(24,16));
ROM(2034) <= std_logic_vector(to_signed(22,16));
ROM(2035) <= std_logic_vector(to_signed(20,16));
ROM(2036) <= std_logic_vector(to_signed(19,16));
ROM(2037) <= std_logic_vector(to_signed(17,16));
ROM(2038) <= std_logic_vector(to_signed(16,16));
ROM(2039) <= std_logic_vector(to_signed(14,16));
ROM(2040) <= std_logic_vector(to_signed(13,16));
ROM(2041) <= std_logic_vector(to_signed(11,16));
ROM(2042) <= std_logic_vector(to_signed(9,16));
ROM(2043) <= std_logic_vector(to_signed(8,16));
ROM(2044) <= std_logic_vector(to_signed(6,16));
ROM(2045) <= std_logic_vector(to_signed(5,16));
ROM(2046) <= std_logic_vector(to_signed(3,16));
ROM(2047) <= std_logic_vector(to_signed(2,16));
ROM(2048) <= std_logic_vector(to_signed(0,16));
ROM(2049) <= std_logic_vector(to_signed(-2,16));
ROM(2050) <= std_logic_vector(to_signed(-3,16));
ROM(2051) <= std_logic_vector(to_signed(-5,16));
ROM(2052) <= std_logic_vector(to_signed(-6,16));
ROM(2053) <= std_logic_vector(to_signed(-8,16));
ROM(2054) <= std_logic_vector(to_signed(-9,16));
ROM(2055) <= std_logic_vector(to_signed(-11,16));
ROM(2056) <= std_logic_vector(to_signed(-13,16));
ROM(2057) <= std_logic_vector(to_signed(-14,16));
ROM(2058) <= std_logic_vector(to_signed(-16,16));
ROM(2059) <= std_logic_vector(to_signed(-17,16));
ROM(2060) <= std_logic_vector(to_signed(-19,16));
ROM(2061) <= std_logic_vector(to_signed(-20,16));
ROM(2062) <= std_logic_vector(to_signed(-22,16));
ROM(2063) <= std_logic_vector(to_signed(-24,16));
ROM(2064) <= std_logic_vector(to_signed(-25,16));
ROM(2065) <= std_logic_vector(to_signed(-27,16));
ROM(2066) <= std_logic_vector(to_signed(-28,16));
ROM(2067) <= std_logic_vector(to_signed(-30,16));
ROM(2068) <= std_logic_vector(to_signed(-31,16));
ROM(2069) <= std_logic_vector(to_signed(-33,16));
ROM(2070) <= std_logic_vector(to_signed(-35,16));
ROM(2071) <= std_logic_vector(to_signed(-36,16));
ROM(2072) <= std_logic_vector(to_signed(-38,16));
ROM(2073) <= std_logic_vector(to_signed(-39,16));
ROM(2074) <= std_logic_vector(to_signed(-41,16));
ROM(2075) <= std_logic_vector(to_signed(-42,16));
ROM(2076) <= std_logic_vector(to_signed(-44,16));
ROM(2077) <= std_logic_vector(to_signed(-46,16));
ROM(2078) <= std_logic_vector(to_signed(-47,16));
ROM(2079) <= std_logic_vector(to_signed(-49,16));
ROM(2080) <= std_logic_vector(to_signed(-50,16));
ROM(2081) <= std_logic_vector(to_signed(-52,16));
ROM(2082) <= std_logic_vector(to_signed(-53,16));
ROM(2083) <= std_logic_vector(to_signed(-55,16));
ROM(2084) <= std_logic_vector(to_signed(-57,16));
ROM(2085) <= std_logic_vector(to_signed(-58,16));
ROM(2086) <= std_logic_vector(to_signed(-60,16));
ROM(2087) <= std_logic_vector(to_signed(-61,16));
ROM(2088) <= std_logic_vector(to_signed(-63,16));
ROM(2089) <= std_logic_vector(to_signed(-64,16));
ROM(2090) <= std_logic_vector(to_signed(-66,16));
ROM(2091) <= std_logic_vector(to_signed(-67,16));
ROM(2092) <= std_logic_vector(to_signed(-69,16));
ROM(2093) <= std_logic_vector(to_signed(-71,16));
ROM(2094) <= std_logic_vector(to_signed(-72,16));
ROM(2095) <= std_logic_vector(to_signed(-74,16));
ROM(2096) <= std_logic_vector(to_signed(-75,16));
ROM(2097) <= std_logic_vector(to_signed(-77,16));
ROM(2098) <= std_logic_vector(to_signed(-78,16));
ROM(2099) <= std_logic_vector(to_signed(-80,16));
ROM(2100) <= std_logic_vector(to_signed(-82,16));
ROM(2101) <= std_logic_vector(to_signed(-83,16));
ROM(2102) <= std_logic_vector(to_signed(-85,16));
ROM(2103) <= std_logic_vector(to_signed(-86,16));
ROM(2104) <= std_logic_vector(to_signed(-88,16));
ROM(2105) <= std_logic_vector(to_signed(-89,16));
ROM(2106) <= std_logic_vector(to_signed(-91,16));
ROM(2107) <= std_logic_vector(to_signed(-93,16));
ROM(2108) <= std_logic_vector(to_signed(-94,16));
ROM(2109) <= std_logic_vector(to_signed(-96,16));
ROM(2110) <= std_logic_vector(to_signed(-97,16));
ROM(2111) <= std_logic_vector(to_signed(-99,16));
ROM(2112) <= std_logic_vector(to_signed(-100,16));
ROM(2113) <= std_logic_vector(to_signed(-102,16));
ROM(2114) <= std_logic_vector(to_signed(-103,16));
ROM(2115) <= std_logic_vector(to_signed(-105,16));
ROM(2116) <= std_logic_vector(to_signed(-107,16));
ROM(2117) <= std_logic_vector(to_signed(-108,16));
ROM(2118) <= std_logic_vector(to_signed(-110,16));
ROM(2119) <= std_logic_vector(to_signed(-111,16));
ROM(2120) <= std_logic_vector(to_signed(-113,16));
ROM(2121) <= std_logic_vector(to_signed(-114,16));
ROM(2122) <= std_logic_vector(to_signed(-116,16));
ROM(2123) <= std_logic_vector(to_signed(-118,16));
ROM(2124) <= std_logic_vector(to_signed(-119,16));
ROM(2125) <= std_logic_vector(to_signed(-121,16));
ROM(2126) <= std_logic_vector(to_signed(-122,16));
ROM(2127) <= std_logic_vector(to_signed(-124,16));
ROM(2128) <= std_logic_vector(to_signed(-125,16));
ROM(2129) <= std_logic_vector(to_signed(-127,16));
ROM(2130) <= std_logic_vector(to_signed(-128,16));
ROM(2131) <= std_logic_vector(to_signed(-130,16));
ROM(2132) <= std_logic_vector(to_signed(-132,16));
ROM(2133) <= std_logic_vector(to_signed(-133,16));
ROM(2134) <= std_logic_vector(to_signed(-135,16));
ROM(2135) <= std_logic_vector(to_signed(-136,16));
ROM(2136) <= std_logic_vector(to_signed(-138,16));
ROM(2137) <= std_logic_vector(to_signed(-139,16));
ROM(2138) <= std_logic_vector(to_signed(-141,16));
ROM(2139) <= std_logic_vector(to_signed(-142,16));
ROM(2140) <= std_logic_vector(to_signed(-144,16));
ROM(2141) <= std_logic_vector(to_signed(-146,16));
ROM(2142) <= std_logic_vector(to_signed(-147,16));
ROM(2143) <= std_logic_vector(to_signed(-149,16));
ROM(2144) <= std_logic_vector(to_signed(-150,16));
ROM(2145) <= std_logic_vector(to_signed(-152,16));
ROM(2146) <= std_logic_vector(to_signed(-153,16));
ROM(2147) <= std_logic_vector(to_signed(-155,16));
ROM(2148) <= std_logic_vector(to_signed(-156,16));
ROM(2149) <= std_logic_vector(to_signed(-158,16));
ROM(2150) <= std_logic_vector(to_signed(-160,16));
ROM(2151) <= std_logic_vector(to_signed(-161,16));
ROM(2152) <= std_logic_vector(to_signed(-163,16));
ROM(2153) <= std_logic_vector(to_signed(-164,16));
ROM(2154) <= std_logic_vector(to_signed(-166,16));
ROM(2155) <= std_logic_vector(to_signed(-167,16));
ROM(2156) <= std_logic_vector(to_signed(-169,16));
ROM(2157) <= std_logic_vector(to_signed(-170,16));
ROM(2158) <= std_logic_vector(to_signed(-172,16));
ROM(2159) <= std_logic_vector(to_signed(-174,16));
ROM(2160) <= std_logic_vector(to_signed(-175,16));
ROM(2161) <= std_logic_vector(to_signed(-177,16));
ROM(2162) <= std_logic_vector(to_signed(-178,16));
ROM(2163) <= std_logic_vector(to_signed(-180,16));
ROM(2164) <= std_logic_vector(to_signed(-181,16));
ROM(2165) <= std_logic_vector(to_signed(-183,16));
ROM(2166) <= std_logic_vector(to_signed(-184,16));
ROM(2167) <= std_logic_vector(to_signed(-186,16));
ROM(2168) <= std_logic_vector(to_signed(-187,16));
ROM(2169) <= std_logic_vector(to_signed(-189,16));
ROM(2170) <= std_logic_vector(to_signed(-191,16));
ROM(2171) <= std_logic_vector(to_signed(-192,16));
ROM(2172) <= std_logic_vector(to_signed(-194,16));
ROM(2173) <= std_logic_vector(to_signed(-195,16));
ROM(2174) <= std_logic_vector(to_signed(-197,16));
ROM(2175) <= std_logic_vector(to_signed(-198,16));
ROM(2176) <= std_logic_vector(to_signed(-200,16));
ROM(2177) <= std_logic_vector(to_signed(-201,16));
ROM(2178) <= std_logic_vector(to_signed(-203,16));
ROM(2179) <= std_logic_vector(to_signed(-204,16));
ROM(2180) <= std_logic_vector(to_signed(-206,16));
ROM(2181) <= std_logic_vector(to_signed(-207,16));
ROM(2182) <= std_logic_vector(to_signed(-209,16));
ROM(2183) <= std_logic_vector(to_signed(-211,16));
ROM(2184) <= std_logic_vector(to_signed(-212,16));
ROM(2185) <= std_logic_vector(to_signed(-214,16));
ROM(2186) <= std_logic_vector(to_signed(-215,16));
ROM(2187) <= std_logic_vector(to_signed(-217,16));
ROM(2188) <= std_logic_vector(to_signed(-218,16));
ROM(2189) <= std_logic_vector(to_signed(-220,16));
ROM(2190) <= std_logic_vector(to_signed(-221,16));
ROM(2191) <= std_logic_vector(to_signed(-223,16));
ROM(2192) <= std_logic_vector(to_signed(-224,16));
ROM(2193) <= std_logic_vector(to_signed(-226,16));
ROM(2194) <= std_logic_vector(to_signed(-227,16));
ROM(2195) <= std_logic_vector(to_signed(-229,16));
ROM(2196) <= std_logic_vector(to_signed(-230,16));
ROM(2197) <= std_logic_vector(to_signed(-232,16));
ROM(2198) <= std_logic_vector(to_signed(-234,16));
ROM(2199) <= std_logic_vector(to_signed(-235,16));
ROM(2200) <= std_logic_vector(to_signed(-237,16));
ROM(2201) <= std_logic_vector(to_signed(-238,16));
ROM(2202) <= std_logic_vector(to_signed(-240,16));
ROM(2203) <= std_logic_vector(to_signed(-241,16));
ROM(2204) <= std_logic_vector(to_signed(-243,16));
ROM(2205) <= std_logic_vector(to_signed(-244,16));
ROM(2206) <= std_logic_vector(to_signed(-246,16));
ROM(2207) <= std_logic_vector(to_signed(-247,16));
ROM(2208) <= std_logic_vector(to_signed(-249,16));
ROM(2209) <= std_logic_vector(to_signed(-250,16));
ROM(2210) <= std_logic_vector(to_signed(-252,16));
ROM(2211) <= std_logic_vector(to_signed(-253,16));
ROM(2212) <= std_logic_vector(to_signed(-255,16));
ROM(2213) <= std_logic_vector(to_signed(-256,16));
ROM(2214) <= std_logic_vector(to_signed(-258,16));
ROM(2215) <= std_logic_vector(to_signed(-259,16));
ROM(2216) <= std_logic_vector(to_signed(-261,16));
ROM(2217) <= std_logic_vector(to_signed(-263,16));
ROM(2218) <= std_logic_vector(to_signed(-264,16));
ROM(2219) <= std_logic_vector(to_signed(-266,16));
ROM(2220) <= std_logic_vector(to_signed(-267,16));
ROM(2221) <= std_logic_vector(to_signed(-269,16));
ROM(2222) <= std_logic_vector(to_signed(-270,16));
ROM(2223) <= std_logic_vector(to_signed(-272,16));
ROM(2224) <= std_logic_vector(to_signed(-273,16));
ROM(2225) <= std_logic_vector(to_signed(-275,16));
ROM(2226) <= std_logic_vector(to_signed(-276,16));
ROM(2227) <= std_logic_vector(to_signed(-278,16));
ROM(2228) <= std_logic_vector(to_signed(-279,16));
ROM(2229) <= std_logic_vector(to_signed(-281,16));
ROM(2230) <= std_logic_vector(to_signed(-282,16));
ROM(2231) <= std_logic_vector(to_signed(-284,16));
ROM(2232) <= std_logic_vector(to_signed(-285,16));
ROM(2233) <= std_logic_vector(to_signed(-287,16));
ROM(2234) <= std_logic_vector(to_signed(-288,16));
ROM(2235) <= std_logic_vector(to_signed(-290,16));
ROM(2236) <= std_logic_vector(to_signed(-291,16));
ROM(2237) <= std_logic_vector(to_signed(-293,16));
ROM(2238) <= std_logic_vector(to_signed(-294,16));
ROM(2239) <= std_logic_vector(to_signed(-296,16));
ROM(2240) <= std_logic_vector(to_signed(-297,16));
ROM(2241) <= std_logic_vector(to_signed(-299,16));
ROM(2242) <= std_logic_vector(to_signed(-300,16));
ROM(2243) <= std_logic_vector(to_signed(-302,16));
ROM(2244) <= std_logic_vector(to_signed(-303,16));
ROM(2245) <= std_logic_vector(to_signed(-305,16));
ROM(2246) <= std_logic_vector(to_signed(-306,16));
ROM(2247) <= std_logic_vector(to_signed(-308,16));
ROM(2248) <= std_logic_vector(to_signed(-309,16));
ROM(2249) <= std_logic_vector(to_signed(-311,16));
ROM(2250) <= std_logic_vector(to_signed(-312,16));
ROM(2251) <= std_logic_vector(to_signed(-314,16));
ROM(2252) <= std_logic_vector(to_signed(-315,16));
ROM(2253) <= std_logic_vector(to_signed(-317,16));
ROM(2254) <= std_logic_vector(to_signed(-318,16));
ROM(2255) <= std_logic_vector(to_signed(-320,16));
ROM(2256) <= std_logic_vector(to_signed(-321,16));
ROM(2257) <= std_logic_vector(to_signed(-323,16));
ROM(2258) <= std_logic_vector(to_signed(-324,16));
ROM(2259) <= std_logic_vector(to_signed(-326,16));
ROM(2260) <= std_logic_vector(to_signed(-327,16));
ROM(2261) <= std_logic_vector(to_signed(-329,16));
ROM(2262) <= std_logic_vector(to_signed(-330,16));
ROM(2263) <= std_logic_vector(to_signed(-332,16));
ROM(2264) <= std_logic_vector(to_signed(-333,16));
ROM(2265) <= std_logic_vector(to_signed(-335,16));
ROM(2266) <= std_logic_vector(to_signed(-336,16));
ROM(2267) <= std_logic_vector(to_signed(-338,16));
ROM(2268) <= std_logic_vector(to_signed(-339,16));
ROM(2269) <= std_logic_vector(to_signed(-341,16));
ROM(2270) <= std_logic_vector(to_signed(-342,16));
ROM(2271) <= std_logic_vector(to_signed(-343,16));
ROM(2272) <= std_logic_vector(to_signed(-345,16));
ROM(2273) <= std_logic_vector(to_signed(-346,16));
ROM(2274) <= std_logic_vector(to_signed(-348,16));
ROM(2275) <= std_logic_vector(to_signed(-349,16));
ROM(2276) <= std_logic_vector(to_signed(-351,16));
ROM(2277) <= std_logic_vector(to_signed(-352,16));
ROM(2278) <= std_logic_vector(to_signed(-354,16));
ROM(2279) <= std_logic_vector(to_signed(-355,16));
ROM(2280) <= std_logic_vector(to_signed(-357,16));
ROM(2281) <= std_logic_vector(to_signed(-358,16));
ROM(2282) <= std_logic_vector(to_signed(-360,16));
ROM(2283) <= std_logic_vector(to_signed(-361,16));
ROM(2284) <= std_logic_vector(to_signed(-363,16));
ROM(2285) <= std_logic_vector(to_signed(-364,16));
ROM(2286) <= std_logic_vector(to_signed(-366,16));
ROM(2287) <= std_logic_vector(to_signed(-367,16));
ROM(2288) <= std_logic_vector(to_signed(-369,16));
ROM(2289) <= std_logic_vector(to_signed(-370,16));
ROM(2290) <= std_logic_vector(to_signed(-371,16));
ROM(2291) <= std_logic_vector(to_signed(-373,16));
ROM(2292) <= std_logic_vector(to_signed(-374,16));
ROM(2293) <= std_logic_vector(to_signed(-376,16));
ROM(2294) <= std_logic_vector(to_signed(-377,16));
ROM(2295) <= std_logic_vector(to_signed(-379,16));
ROM(2296) <= std_logic_vector(to_signed(-380,16));
ROM(2297) <= std_logic_vector(to_signed(-382,16));
ROM(2298) <= std_logic_vector(to_signed(-383,16));
ROM(2299) <= std_logic_vector(to_signed(-385,16));
ROM(2300) <= std_logic_vector(to_signed(-386,16));
ROM(2301) <= std_logic_vector(to_signed(-388,16));
ROM(2302) <= std_logic_vector(to_signed(-389,16));
ROM(2303) <= std_logic_vector(to_signed(-390,16));
ROM(2304) <= std_logic_vector(to_signed(-392,16));
ROM(2305) <= std_logic_vector(to_signed(-393,16));
ROM(2306) <= std_logic_vector(to_signed(-395,16));
ROM(2307) <= std_logic_vector(to_signed(-396,16));
ROM(2308) <= std_logic_vector(to_signed(-398,16));
ROM(2309) <= std_logic_vector(to_signed(-399,16));
ROM(2310) <= std_logic_vector(to_signed(-401,16));
ROM(2311) <= std_logic_vector(to_signed(-402,16));
ROM(2312) <= std_logic_vector(to_signed(-403,16));
ROM(2313) <= std_logic_vector(to_signed(-405,16));
ROM(2314) <= std_logic_vector(to_signed(-406,16));
ROM(2315) <= std_logic_vector(to_signed(-408,16));
ROM(2316) <= std_logic_vector(to_signed(-409,16));
ROM(2317) <= std_logic_vector(to_signed(-411,16));
ROM(2318) <= std_logic_vector(to_signed(-412,16));
ROM(2319) <= std_logic_vector(to_signed(-414,16));
ROM(2320) <= std_logic_vector(to_signed(-415,16));
ROM(2321) <= std_logic_vector(to_signed(-416,16));
ROM(2322) <= std_logic_vector(to_signed(-418,16));
ROM(2323) <= std_logic_vector(to_signed(-419,16));
ROM(2324) <= std_logic_vector(to_signed(-421,16));
ROM(2325) <= std_logic_vector(to_signed(-422,16));
ROM(2326) <= std_logic_vector(to_signed(-424,16));
ROM(2327) <= std_logic_vector(to_signed(-425,16));
ROM(2328) <= std_logic_vector(to_signed(-426,16));
ROM(2329) <= std_logic_vector(to_signed(-428,16));
ROM(2330) <= std_logic_vector(to_signed(-429,16));
ROM(2331) <= std_logic_vector(to_signed(-431,16));
ROM(2332) <= std_logic_vector(to_signed(-432,16));
ROM(2333) <= std_logic_vector(to_signed(-434,16));
ROM(2334) <= std_logic_vector(to_signed(-435,16));
ROM(2335) <= std_logic_vector(to_signed(-436,16));
ROM(2336) <= std_logic_vector(to_signed(-438,16));
ROM(2337) <= std_logic_vector(to_signed(-439,16));
ROM(2338) <= std_logic_vector(to_signed(-441,16));
ROM(2339) <= std_logic_vector(to_signed(-442,16));
ROM(2340) <= std_logic_vector(to_signed(-443,16));
ROM(2341) <= std_logic_vector(to_signed(-445,16));
ROM(2342) <= std_logic_vector(to_signed(-446,16));
ROM(2343) <= std_logic_vector(to_signed(-448,16));
ROM(2344) <= std_logic_vector(to_signed(-449,16));
ROM(2345) <= std_logic_vector(to_signed(-451,16));
ROM(2346) <= std_logic_vector(to_signed(-452,16));
ROM(2347) <= std_logic_vector(to_signed(-453,16));
ROM(2348) <= std_logic_vector(to_signed(-455,16));
ROM(2349) <= std_logic_vector(to_signed(-456,16));
ROM(2350) <= std_logic_vector(to_signed(-458,16));
ROM(2351) <= std_logic_vector(to_signed(-459,16));
ROM(2352) <= std_logic_vector(to_signed(-460,16));
ROM(2353) <= std_logic_vector(to_signed(-462,16));
ROM(2354) <= std_logic_vector(to_signed(-463,16));
ROM(2355) <= std_logic_vector(to_signed(-465,16));
ROM(2356) <= std_logic_vector(to_signed(-466,16));
ROM(2357) <= std_logic_vector(to_signed(-467,16));
ROM(2358) <= std_logic_vector(to_signed(-469,16));
ROM(2359) <= std_logic_vector(to_signed(-470,16));
ROM(2360) <= std_logic_vector(to_signed(-472,16));
ROM(2361) <= std_logic_vector(to_signed(-473,16));
ROM(2362) <= std_logic_vector(to_signed(-474,16));
ROM(2363) <= std_logic_vector(to_signed(-476,16));
ROM(2364) <= std_logic_vector(to_signed(-477,16));
ROM(2365) <= std_logic_vector(to_signed(-479,16));
ROM(2366) <= std_logic_vector(to_signed(-480,16));
ROM(2367) <= std_logic_vector(to_signed(-481,16));
ROM(2368) <= std_logic_vector(to_signed(-483,16));
ROM(2369) <= std_logic_vector(to_signed(-484,16));
ROM(2370) <= std_logic_vector(to_signed(-485,16));
ROM(2371) <= std_logic_vector(to_signed(-487,16));
ROM(2372) <= std_logic_vector(to_signed(-488,16));
ROM(2373) <= std_logic_vector(to_signed(-490,16));
ROM(2374) <= std_logic_vector(to_signed(-491,16));
ROM(2375) <= std_logic_vector(to_signed(-492,16));
ROM(2376) <= std_logic_vector(to_signed(-494,16));
ROM(2377) <= std_logic_vector(to_signed(-495,16));
ROM(2378) <= std_logic_vector(to_signed(-497,16));
ROM(2379) <= std_logic_vector(to_signed(-498,16));
ROM(2380) <= std_logic_vector(to_signed(-499,16));
ROM(2381) <= std_logic_vector(to_signed(-501,16));
ROM(2382) <= std_logic_vector(to_signed(-502,16));
ROM(2383) <= std_logic_vector(to_signed(-503,16));
ROM(2384) <= std_logic_vector(to_signed(-505,16));
ROM(2385) <= std_logic_vector(to_signed(-506,16));
ROM(2386) <= std_logic_vector(to_signed(-507,16));
ROM(2387) <= std_logic_vector(to_signed(-509,16));
ROM(2388) <= std_logic_vector(to_signed(-510,16));
ROM(2389) <= std_logic_vector(to_signed(-512,16));
ROM(2390) <= std_logic_vector(to_signed(-513,16));
ROM(2391) <= std_logic_vector(to_signed(-514,16));
ROM(2392) <= std_logic_vector(to_signed(-516,16));
ROM(2393) <= std_logic_vector(to_signed(-517,16));
ROM(2394) <= std_logic_vector(to_signed(-518,16));
ROM(2395) <= std_logic_vector(to_signed(-520,16));
ROM(2396) <= std_logic_vector(to_signed(-521,16));
ROM(2397) <= std_logic_vector(to_signed(-522,16));
ROM(2398) <= std_logic_vector(to_signed(-524,16));
ROM(2399) <= std_logic_vector(to_signed(-525,16));
ROM(2400) <= std_logic_vector(to_signed(-526,16));
ROM(2401) <= std_logic_vector(to_signed(-528,16));
ROM(2402) <= std_logic_vector(to_signed(-529,16));
ROM(2403) <= std_logic_vector(to_signed(-530,16));
ROM(2404) <= std_logic_vector(to_signed(-532,16));
ROM(2405) <= std_logic_vector(to_signed(-533,16));
ROM(2406) <= std_logic_vector(to_signed(-535,16));
ROM(2407) <= std_logic_vector(to_signed(-536,16));
ROM(2408) <= std_logic_vector(to_signed(-537,16));
ROM(2409) <= std_logic_vector(to_signed(-539,16));
ROM(2410) <= std_logic_vector(to_signed(-540,16));
ROM(2411) <= std_logic_vector(to_signed(-541,16));
ROM(2412) <= std_logic_vector(to_signed(-543,16));
ROM(2413) <= std_logic_vector(to_signed(-544,16));
ROM(2414) <= std_logic_vector(to_signed(-545,16));
ROM(2415) <= std_logic_vector(to_signed(-547,16));
ROM(2416) <= std_logic_vector(to_signed(-548,16));
ROM(2417) <= std_logic_vector(to_signed(-549,16));
ROM(2418) <= std_logic_vector(to_signed(-550,16));
ROM(2419) <= std_logic_vector(to_signed(-552,16));
ROM(2420) <= std_logic_vector(to_signed(-553,16));
ROM(2421) <= std_logic_vector(to_signed(-554,16));
ROM(2422) <= std_logic_vector(to_signed(-556,16));
ROM(2423) <= std_logic_vector(to_signed(-557,16));
ROM(2424) <= std_logic_vector(to_signed(-558,16));
ROM(2425) <= std_logic_vector(to_signed(-560,16));
ROM(2426) <= std_logic_vector(to_signed(-561,16));
ROM(2427) <= std_logic_vector(to_signed(-562,16));
ROM(2428) <= std_logic_vector(to_signed(-564,16));
ROM(2429) <= std_logic_vector(to_signed(-565,16));
ROM(2430) <= std_logic_vector(to_signed(-566,16));
ROM(2431) <= std_logic_vector(to_signed(-568,16));
ROM(2432) <= std_logic_vector(to_signed(-569,16));
ROM(2433) <= std_logic_vector(to_signed(-570,16));
ROM(2434) <= std_logic_vector(to_signed(-572,16));
ROM(2435) <= std_logic_vector(to_signed(-573,16));
ROM(2436) <= std_logic_vector(to_signed(-574,16));
ROM(2437) <= std_logic_vector(to_signed(-575,16));
ROM(2438) <= std_logic_vector(to_signed(-577,16));
ROM(2439) <= std_logic_vector(to_signed(-578,16));
ROM(2440) <= std_logic_vector(to_signed(-579,16));
ROM(2441) <= std_logic_vector(to_signed(-581,16));
ROM(2442) <= std_logic_vector(to_signed(-582,16));
ROM(2443) <= std_logic_vector(to_signed(-583,16));
ROM(2444) <= std_logic_vector(to_signed(-584,16));
ROM(2445) <= std_logic_vector(to_signed(-586,16));
ROM(2446) <= std_logic_vector(to_signed(-587,16));
ROM(2447) <= std_logic_vector(to_signed(-588,16));
ROM(2448) <= std_logic_vector(to_signed(-590,16));
ROM(2449) <= std_logic_vector(to_signed(-591,16));
ROM(2450) <= std_logic_vector(to_signed(-592,16));
ROM(2451) <= std_logic_vector(to_signed(-593,16));
ROM(2452) <= std_logic_vector(to_signed(-595,16));
ROM(2453) <= std_logic_vector(to_signed(-596,16));
ROM(2454) <= std_logic_vector(to_signed(-597,16));
ROM(2455) <= std_logic_vector(to_signed(-599,16));
ROM(2456) <= std_logic_vector(to_signed(-600,16));
ROM(2457) <= std_logic_vector(to_signed(-601,16));
ROM(2458) <= std_logic_vector(to_signed(-602,16));
ROM(2459) <= std_logic_vector(to_signed(-604,16));
ROM(2460) <= std_logic_vector(to_signed(-605,16));
ROM(2461) <= std_logic_vector(to_signed(-606,16));
ROM(2462) <= std_logic_vector(to_signed(-607,16));
ROM(2463) <= std_logic_vector(to_signed(-609,16));
ROM(2464) <= std_logic_vector(to_signed(-610,16));
ROM(2465) <= std_logic_vector(to_signed(-611,16));
ROM(2466) <= std_logic_vector(to_signed(-613,16));
ROM(2467) <= std_logic_vector(to_signed(-614,16));
ROM(2468) <= std_logic_vector(to_signed(-615,16));
ROM(2469) <= std_logic_vector(to_signed(-616,16));
ROM(2470) <= std_logic_vector(to_signed(-618,16));
ROM(2471) <= std_logic_vector(to_signed(-619,16));
ROM(2472) <= std_logic_vector(to_signed(-620,16));
ROM(2473) <= std_logic_vector(to_signed(-621,16));
ROM(2474) <= std_logic_vector(to_signed(-623,16));
ROM(2475) <= std_logic_vector(to_signed(-624,16));
ROM(2476) <= std_logic_vector(to_signed(-625,16));
ROM(2477) <= std_logic_vector(to_signed(-626,16));
ROM(2478) <= std_logic_vector(to_signed(-628,16));
ROM(2479) <= std_logic_vector(to_signed(-629,16));
ROM(2480) <= std_logic_vector(to_signed(-630,16));
ROM(2481) <= std_logic_vector(to_signed(-631,16));
ROM(2482) <= std_logic_vector(to_signed(-632,16));
ROM(2483) <= std_logic_vector(to_signed(-634,16));
ROM(2484) <= std_logic_vector(to_signed(-635,16));
ROM(2485) <= std_logic_vector(to_signed(-636,16));
ROM(2486) <= std_logic_vector(to_signed(-637,16));
ROM(2487) <= std_logic_vector(to_signed(-639,16));
ROM(2488) <= std_logic_vector(to_signed(-640,16));
ROM(2489) <= std_logic_vector(to_signed(-641,16));
ROM(2490) <= std_logic_vector(to_signed(-642,16));
ROM(2491) <= std_logic_vector(to_signed(-644,16));
ROM(2492) <= std_logic_vector(to_signed(-645,16));
ROM(2493) <= std_logic_vector(to_signed(-646,16));
ROM(2494) <= std_logic_vector(to_signed(-647,16));
ROM(2495) <= std_logic_vector(to_signed(-648,16));
ROM(2496) <= std_logic_vector(to_signed(-650,16));
ROM(2497) <= std_logic_vector(to_signed(-651,16));
ROM(2498) <= std_logic_vector(to_signed(-652,16));
ROM(2499) <= std_logic_vector(to_signed(-653,16));
ROM(2500) <= std_logic_vector(to_signed(-654,16));
ROM(2501) <= std_logic_vector(to_signed(-656,16));
ROM(2502) <= std_logic_vector(to_signed(-657,16));
ROM(2503) <= std_logic_vector(to_signed(-658,16));
ROM(2504) <= std_logic_vector(to_signed(-659,16));
ROM(2505) <= std_logic_vector(to_signed(-660,16));
ROM(2506) <= std_logic_vector(to_signed(-662,16));
ROM(2507) <= std_logic_vector(to_signed(-663,16));
ROM(2508) <= std_logic_vector(to_signed(-664,16));
ROM(2509) <= std_logic_vector(to_signed(-665,16));
ROM(2510) <= std_logic_vector(to_signed(-666,16));
ROM(2511) <= std_logic_vector(to_signed(-668,16));
ROM(2512) <= std_logic_vector(to_signed(-669,16));
ROM(2513) <= std_logic_vector(to_signed(-670,16));
ROM(2514) <= std_logic_vector(to_signed(-671,16));
ROM(2515) <= std_logic_vector(to_signed(-672,16));
ROM(2516) <= std_logic_vector(to_signed(-674,16));
ROM(2517) <= std_logic_vector(to_signed(-675,16));
ROM(2518) <= std_logic_vector(to_signed(-676,16));
ROM(2519) <= std_logic_vector(to_signed(-677,16));
ROM(2520) <= std_logic_vector(to_signed(-678,16));
ROM(2521) <= std_logic_vector(to_signed(-679,16));
ROM(2522) <= std_logic_vector(to_signed(-681,16));
ROM(2523) <= std_logic_vector(to_signed(-682,16));
ROM(2524) <= std_logic_vector(to_signed(-683,16));
ROM(2525) <= std_logic_vector(to_signed(-684,16));
ROM(2526) <= std_logic_vector(to_signed(-685,16));
ROM(2527) <= std_logic_vector(to_signed(-687,16));
ROM(2528) <= std_logic_vector(to_signed(-688,16));
ROM(2529) <= std_logic_vector(to_signed(-689,16));
ROM(2530) <= std_logic_vector(to_signed(-690,16));
ROM(2531) <= std_logic_vector(to_signed(-691,16));
ROM(2532) <= std_logic_vector(to_signed(-692,16));
ROM(2533) <= std_logic_vector(to_signed(-693,16));
ROM(2534) <= std_logic_vector(to_signed(-695,16));
ROM(2535) <= std_logic_vector(to_signed(-696,16));
ROM(2536) <= std_logic_vector(to_signed(-697,16));
ROM(2537) <= std_logic_vector(to_signed(-698,16));
ROM(2538) <= std_logic_vector(to_signed(-699,16));
ROM(2539) <= std_logic_vector(to_signed(-700,16));
ROM(2540) <= std_logic_vector(to_signed(-702,16));
ROM(2541) <= std_logic_vector(to_signed(-703,16));
ROM(2542) <= std_logic_vector(to_signed(-704,16));
ROM(2543) <= std_logic_vector(to_signed(-705,16));
ROM(2544) <= std_logic_vector(to_signed(-706,16));
ROM(2545) <= std_logic_vector(to_signed(-707,16));
ROM(2546) <= std_logic_vector(to_signed(-708,16));
ROM(2547) <= std_logic_vector(to_signed(-709,16));
ROM(2548) <= std_logic_vector(to_signed(-711,16));
ROM(2549) <= std_logic_vector(to_signed(-712,16));
ROM(2550) <= std_logic_vector(to_signed(-713,16));
ROM(2551) <= std_logic_vector(to_signed(-714,16));
ROM(2552) <= std_logic_vector(to_signed(-715,16));
ROM(2553) <= std_logic_vector(to_signed(-716,16));
ROM(2554) <= std_logic_vector(to_signed(-717,16));
ROM(2555) <= std_logic_vector(to_signed(-719,16));
ROM(2556) <= std_logic_vector(to_signed(-720,16));
ROM(2557) <= std_logic_vector(to_signed(-721,16));
ROM(2558) <= std_logic_vector(to_signed(-722,16));
ROM(2559) <= std_logic_vector(to_signed(-723,16));
ROM(2560) <= std_logic_vector(to_signed(-724,16));
ROM(2561) <= std_logic_vector(to_signed(-725,16));
ROM(2562) <= std_logic_vector(to_signed(-726,16));
ROM(2563) <= std_logic_vector(to_signed(-727,16));
ROM(2564) <= std_logic_vector(to_signed(-729,16));
ROM(2565) <= std_logic_vector(to_signed(-730,16));
ROM(2566) <= std_logic_vector(to_signed(-731,16));
ROM(2567) <= std_logic_vector(to_signed(-732,16));
ROM(2568) <= std_logic_vector(to_signed(-733,16));
ROM(2569) <= std_logic_vector(to_signed(-734,16));
ROM(2570) <= std_logic_vector(to_signed(-735,16));
ROM(2571) <= std_logic_vector(to_signed(-736,16));
ROM(2572) <= std_logic_vector(to_signed(-737,16));
ROM(2573) <= std_logic_vector(to_signed(-738,16));
ROM(2574) <= std_logic_vector(to_signed(-739,16));
ROM(2575) <= std_logic_vector(to_signed(-741,16));
ROM(2576) <= std_logic_vector(to_signed(-742,16));
ROM(2577) <= std_logic_vector(to_signed(-743,16));
ROM(2578) <= std_logic_vector(to_signed(-744,16));
ROM(2579) <= std_logic_vector(to_signed(-745,16));
ROM(2580) <= std_logic_vector(to_signed(-746,16));
ROM(2581) <= std_logic_vector(to_signed(-747,16));
ROM(2582) <= std_logic_vector(to_signed(-748,16));
ROM(2583) <= std_logic_vector(to_signed(-749,16));
ROM(2584) <= std_logic_vector(to_signed(-750,16));
ROM(2585) <= std_logic_vector(to_signed(-751,16));
ROM(2586) <= std_logic_vector(to_signed(-752,16));
ROM(2587) <= std_logic_vector(to_signed(-753,16));
ROM(2588) <= std_logic_vector(to_signed(-755,16));
ROM(2589) <= std_logic_vector(to_signed(-756,16));
ROM(2590) <= std_logic_vector(to_signed(-757,16));
ROM(2591) <= std_logic_vector(to_signed(-758,16));
ROM(2592) <= std_logic_vector(to_signed(-759,16));
ROM(2593) <= std_logic_vector(to_signed(-760,16));
ROM(2594) <= std_logic_vector(to_signed(-761,16));
ROM(2595) <= std_logic_vector(to_signed(-762,16));
ROM(2596) <= std_logic_vector(to_signed(-763,16));
ROM(2597) <= std_logic_vector(to_signed(-764,16));
ROM(2598) <= std_logic_vector(to_signed(-765,16));
ROM(2599) <= std_logic_vector(to_signed(-766,16));
ROM(2600) <= std_logic_vector(to_signed(-767,16));
ROM(2601) <= std_logic_vector(to_signed(-768,16));
ROM(2602) <= std_logic_vector(to_signed(-769,16));
ROM(2603) <= std_logic_vector(to_signed(-770,16));
ROM(2604) <= std_logic_vector(to_signed(-771,16));
ROM(2605) <= std_logic_vector(to_signed(-772,16));
ROM(2606) <= std_logic_vector(to_signed(-773,16));
ROM(2607) <= std_logic_vector(to_signed(-774,16));
ROM(2608) <= std_logic_vector(to_signed(-775,16));
ROM(2609) <= std_logic_vector(to_signed(-776,16));
ROM(2610) <= std_logic_vector(to_signed(-777,16));
ROM(2611) <= std_logic_vector(to_signed(-778,16));
ROM(2612) <= std_logic_vector(to_signed(-779,16));
ROM(2613) <= std_logic_vector(to_signed(-780,16));
ROM(2614) <= std_logic_vector(to_signed(-782,16));
ROM(2615) <= std_logic_vector(to_signed(-783,16));
ROM(2616) <= std_logic_vector(to_signed(-784,16));
ROM(2617) <= std_logic_vector(to_signed(-785,16));
ROM(2618) <= std_logic_vector(to_signed(-786,16));
ROM(2619) <= std_logic_vector(to_signed(-787,16));
ROM(2620) <= std_logic_vector(to_signed(-788,16));
ROM(2621) <= std_logic_vector(to_signed(-789,16));
ROM(2622) <= std_logic_vector(to_signed(-790,16));
ROM(2623) <= std_logic_vector(to_signed(-791,16));
ROM(2624) <= std_logic_vector(to_signed(-792,16));
ROM(2625) <= std_logic_vector(to_signed(-793,16));
ROM(2626) <= std_logic_vector(to_signed(-794,16));
ROM(2627) <= std_logic_vector(to_signed(-795,16));
ROM(2628) <= std_logic_vector(to_signed(-796,16));
ROM(2629) <= std_logic_vector(to_signed(-797,16));
ROM(2630) <= std_logic_vector(to_signed(-798,16));
ROM(2631) <= std_logic_vector(to_signed(-798,16));
ROM(2632) <= std_logic_vector(to_signed(-799,16));
ROM(2633) <= std_logic_vector(to_signed(-800,16));
ROM(2634) <= std_logic_vector(to_signed(-801,16));
ROM(2635) <= std_logic_vector(to_signed(-802,16));
ROM(2636) <= std_logic_vector(to_signed(-803,16));
ROM(2637) <= std_logic_vector(to_signed(-804,16));
ROM(2638) <= std_logic_vector(to_signed(-805,16));
ROM(2639) <= std_logic_vector(to_signed(-806,16));
ROM(2640) <= std_logic_vector(to_signed(-807,16));
ROM(2641) <= std_logic_vector(to_signed(-808,16));
ROM(2642) <= std_logic_vector(to_signed(-809,16));
ROM(2643) <= std_logic_vector(to_signed(-810,16));
ROM(2644) <= std_logic_vector(to_signed(-811,16));
ROM(2645) <= std_logic_vector(to_signed(-812,16));
ROM(2646) <= std_logic_vector(to_signed(-813,16));
ROM(2647) <= std_logic_vector(to_signed(-814,16));
ROM(2648) <= std_logic_vector(to_signed(-815,16));
ROM(2649) <= std_logic_vector(to_signed(-816,16));
ROM(2650) <= std_logic_vector(to_signed(-817,16));
ROM(2651) <= std_logic_vector(to_signed(-818,16));
ROM(2652) <= std_logic_vector(to_signed(-819,16));
ROM(2653) <= std_logic_vector(to_signed(-820,16));
ROM(2654) <= std_logic_vector(to_signed(-821,16));
ROM(2655) <= std_logic_vector(to_signed(-822,16));
ROM(2656) <= std_logic_vector(to_signed(-822,16));
ROM(2657) <= std_logic_vector(to_signed(-823,16));
ROM(2658) <= std_logic_vector(to_signed(-824,16));
ROM(2659) <= std_logic_vector(to_signed(-825,16));
ROM(2660) <= std_logic_vector(to_signed(-826,16));
ROM(2661) <= std_logic_vector(to_signed(-827,16));
ROM(2662) <= std_logic_vector(to_signed(-828,16));
ROM(2663) <= std_logic_vector(to_signed(-829,16));
ROM(2664) <= std_logic_vector(to_signed(-830,16));
ROM(2665) <= std_logic_vector(to_signed(-831,16));
ROM(2666) <= std_logic_vector(to_signed(-832,16));
ROM(2667) <= std_logic_vector(to_signed(-833,16));
ROM(2668) <= std_logic_vector(to_signed(-834,16));
ROM(2669) <= std_logic_vector(to_signed(-834,16));
ROM(2670) <= std_logic_vector(to_signed(-835,16));
ROM(2671) <= std_logic_vector(to_signed(-836,16));
ROM(2672) <= std_logic_vector(to_signed(-837,16));
ROM(2673) <= std_logic_vector(to_signed(-838,16));
ROM(2674) <= std_logic_vector(to_signed(-839,16));
ROM(2675) <= std_logic_vector(to_signed(-840,16));
ROM(2676) <= std_logic_vector(to_signed(-841,16));
ROM(2677) <= std_logic_vector(to_signed(-842,16));
ROM(2678) <= std_logic_vector(to_signed(-843,16));
ROM(2679) <= std_logic_vector(to_signed(-843,16));
ROM(2680) <= std_logic_vector(to_signed(-844,16));
ROM(2681) <= std_logic_vector(to_signed(-845,16));
ROM(2682) <= std_logic_vector(to_signed(-846,16));
ROM(2683) <= std_logic_vector(to_signed(-847,16));
ROM(2684) <= std_logic_vector(to_signed(-848,16));
ROM(2685) <= std_logic_vector(to_signed(-849,16));
ROM(2686) <= std_logic_vector(to_signed(-850,16));
ROM(2687) <= std_logic_vector(to_signed(-851,16));
ROM(2688) <= std_logic_vector(to_signed(-851,16));
ROM(2689) <= std_logic_vector(to_signed(-852,16));
ROM(2690) <= std_logic_vector(to_signed(-853,16));
ROM(2691) <= std_logic_vector(to_signed(-854,16));
ROM(2692) <= std_logic_vector(to_signed(-855,16));
ROM(2693) <= std_logic_vector(to_signed(-856,16));
ROM(2694) <= std_logic_vector(to_signed(-857,16));
ROM(2695) <= std_logic_vector(to_signed(-857,16));
ROM(2696) <= std_logic_vector(to_signed(-858,16));
ROM(2697) <= std_logic_vector(to_signed(-859,16));
ROM(2698) <= std_logic_vector(to_signed(-860,16));
ROM(2699) <= std_logic_vector(to_signed(-861,16));
ROM(2700) <= std_logic_vector(to_signed(-862,16));
ROM(2701) <= std_logic_vector(to_signed(-863,16));
ROM(2702) <= std_logic_vector(to_signed(-863,16));
ROM(2703) <= std_logic_vector(to_signed(-864,16));
ROM(2704) <= std_logic_vector(to_signed(-865,16));
ROM(2705) <= std_logic_vector(to_signed(-866,16));
ROM(2706) <= std_logic_vector(to_signed(-867,16));
ROM(2707) <= std_logic_vector(to_signed(-868,16));
ROM(2708) <= std_logic_vector(to_signed(-868,16));
ROM(2709) <= std_logic_vector(to_signed(-869,16));
ROM(2710) <= std_logic_vector(to_signed(-870,16));
ROM(2711) <= std_logic_vector(to_signed(-871,16));
ROM(2712) <= std_logic_vector(to_signed(-872,16));
ROM(2713) <= std_logic_vector(to_signed(-873,16));
ROM(2714) <= std_logic_vector(to_signed(-873,16));
ROM(2715) <= std_logic_vector(to_signed(-874,16));
ROM(2716) <= std_logic_vector(to_signed(-875,16));
ROM(2717) <= std_logic_vector(to_signed(-876,16));
ROM(2718) <= std_logic_vector(to_signed(-877,16));
ROM(2719) <= std_logic_vector(to_signed(-878,16));
ROM(2720) <= std_logic_vector(to_signed(-878,16));
ROM(2721) <= std_logic_vector(to_signed(-879,16));
ROM(2722) <= std_logic_vector(to_signed(-880,16));
ROM(2723) <= std_logic_vector(to_signed(-881,16));
ROM(2724) <= std_logic_vector(to_signed(-882,16));
ROM(2725) <= std_logic_vector(to_signed(-882,16));
ROM(2726) <= std_logic_vector(to_signed(-883,16));
ROM(2727) <= std_logic_vector(to_signed(-884,16));
ROM(2728) <= std_logic_vector(to_signed(-885,16));
ROM(2729) <= std_logic_vector(to_signed(-885,16));
ROM(2730) <= std_logic_vector(to_signed(-886,16));
ROM(2731) <= std_logic_vector(to_signed(-887,16));
ROM(2732) <= std_logic_vector(to_signed(-888,16));
ROM(2733) <= std_logic_vector(to_signed(-889,16));
ROM(2734) <= std_logic_vector(to_signed(-889,16));
ROM(2735) <= std_logic_vector(to_signed(-890,16));
ROM(2736) <= std_logic_vector(to_signed(-891,16));
ROM(2737) <= std_logic_vector(to_signed(-892,16));
ROM(2738) <= std_logic_vector(to_signed(-893,16));
ROM(2739) <= std_logic_vector(to_signed(-893,16));
ROM(2740) <= std_logic_vector(to_signed(-894,16));
ROM(2741) <= std_logic_vector(to_signed(-895,16));
ROM(2742) <= std_logic_vector(to_signed(-896,16));
ROM(2743) <= std_logic_vector(to_signed(-896,16));
ROM(2744) <= std_logic_vector(to_signed(-897,16));
ROM(2745) <= std_logic_vector(to_signed(-898,16));
ROM(2746) <= std_logic_vector(to_signed(-899,16));
ROM(2747) <= std_logic_vector(to_signed(-899,16));
ROM(2748) <= std_logic_vector(to_signed(-900,16));
ROM(2749) <= std_logic_vector(to_signed(-901,16));
ROM(2750) <= std_logic_vector(to_signed(-902,16));
ROM(2751) <= std_logic_vector(to_signed(-902,16));
ROM(2752) <= std_logic_vector(to_signed(-903,16));
ROM(2753) <= std_logic_vector(to_signed(-904,16));
ROM(2754) <= std_logic_vector(to_signed(-905,16));
ROM(2755) <= std_logic_vector(to_signed(-905,16));
ROM(2756) <= std_logic_vector(to_signed(-906,16));
ROM(2757) <= std_logic_vector(to_signed(-907,16));
ROM(2758) <= std_logic_vector(to_signed(-907,16));
ROM(2759) <= std_logic_vector(to_signed(-908,16));
ROM(2760) <= std_logic_vector(to_signed(-909,16));
ROM(2761) <= std_logic_vector(to_signed(-910,16));
ROM(2762) <= std_logic_vector(to_signed(-910,16));
ROM(2763) <= std_logic_vector(to_signed(-911,16));
ROM(2764) <= std_logic_vector(to_signed(-912,16));
ROM(2765) <= std_logic_vector(to_signed(-913,16));
ROM(2766) <= std_logic_vector(to_signed(-913,16));
ROM(2767) <= std_logic_vector(to_signed(-914,16));
ROM(2768) <= std_logic_vector(to_signed(-915,16));
ROM(2769) <= std_logic_vector(to_signed(-915,16));
ROM(2770) <= std_logic_vector(to_signed(-916,16));
ROM(2771) <= std_logic_vector(to_signed(-917,16));
ROM(2772) <= std_logic_vector(to_signed(-917,16));
ROM(2773) <= std_logic_vector(to_signed(-918,16));
ROM(2774) <= std_logic_vector(to_signed(-919,16));
ROM(2775) <= std_logic_vector(to_signed(-920,16));
ROM(2776) <= std_logic_vector(to_signed(-920,16));
ROM(2777) <= std_logic_vector(to_signed(-921,16));
ROM(2778) <= std_logic_vector(to_signed(-922,16));
ROM(2779) <= std_logic_vector(to_signed(-922,16));
ROM(2780) <= std_logic_vector(to_signed(-923,16));
ROM(2781) <= std_logic_vector(to_signed(-924,16));
ROM(2782) <= std_logic_vector(to_signed(-924,16));
ROM(2783) <= std_logic_vector(to_signed(-925,16));
ROM(2784) <= std_logic_vector(to_signed(-926,16));
ROM(2785) <= std_logic_vector(to_signed(-926,16));
ROM(2786) <= std_logic_vector(to_signed(-927,16));
ROM(2787) <= std_logic_vector(to_signed(-928,16));
ROM(2788) <= std_logic_vector(to_signed(-928,16));
ROM(2789) <= std_logic_vector(to_signed(-929,16));
ROM(2790) <= std_logic_vector(to_signed(-930,16));
ROM(2791) <= std_logic_vector(to_signed(-930,16));
ROM(2792) <= std_logic_vector(to_signed(-931,16));
ROM(2793) <= std_logic_vector(to_signed(-932,16));
ROM(2794) <= std_logic_vector(to_signed(-932,16));
ROM(2795) <= std_logic_vector(to_signed(-933,16));
ROM(2796) <= std_logic_vector(to_signed(-934,16));
ROM(2797) <= std_logic_vector(to_signed(-934,16));
ROM(2798) <= std_logic_vector(to_signed(-935,16));
ROM(2799) <= std_logic_vector(to_signed(-936,16));
ROM(2800) <= std_logic_vector(to_signed(-936,16));
ROM(2801) <= std_logic_vector(to_signed(-937,16));
ROM(2802) <= std_logic_vector(to_signed(-937,16));
ROM(2803) <= std_logic_vector(to_signed(-938,16));
ROM(2804) <= std_logic_vector(to_signed(-939,16));
ROM(2805) <= std_logic_vector(to_signed(-939,16));
ROM(2806) <= std_logic_vector(to_signed(-940,16));
ROM(2807) <= std_logic_vector(to_signed(-941,16));
ROM(2808) <= std_logic_vector(to_signed(-941,16));
ROM(2809) <= std_logic_vector(to_signed(-942,16));
ROM(2810) <= std_logic_vector(to_signed(-942,16));
ROM(2811) <= std_logic_vector(to_signed(-943,16));
ROM(2812) <= std_logic_vector(to_signed(-944,16));
ROM(2813) <= std_logic_vector(to_signed(-944,16));
ROM(2814) <= std_logic_vector(to_signed(-945,16));
ROM(2815) <= std_logic_vector(to_signed(-945,16));
ROM(2816) <= std_logic_vector(to_signed(-946,16));
ROM(2817) <= std_logic_vector(to_signed(-947,16));
ROM(2818) <= std_logic_vector(to_signed(-947,16));
ROM(2819) <= std_logic_vector(to_signed(-948,16));
ROM(2820) <= std_logic_vector(to_signed(-948,16));
ROM(2821) <= std_logic_vector(to_signed(-949,16));
ROM(2822) <= std_logic_vector(to_signed(-950,16));
ROM(2823) <= std_logic_vector(to_signed(-950,16));
ROM(2824) <= std_logic_vector(to_signed(-951,16));
ROM(2825) <= std_logic_vector(to_signed(-951,16));
ROM(2826) <= std_logic_vector(to_signed(-952,16));
ROM(2827) <= std_logic_vector(to_signed(-953,16));
ROM(2828) <= std_logic_vector(to_signed(-953,16));
ROM(2829) <= std_logic_vector(to_signed(-954,16));
ROM(2830) <= std_logic_vector(to_signed(-954,16));
ROM(2831) <= std_logic_vector(to_signed(-955,16));
ROM(2832) <= std_logic_vector(to_signed(-955,16));
ROM(2833) <= std_logic_vector(to_signed(-956,16));
ROM(2834) <= std_logic_vector(to_signed(-957,16));
ROM(2835) <= std_logic_vector(to_signed(-957,16));
ROM(2836) <= std_logic_vector(to_signed(-958,16));
ROM(2837) <= std_logic_vector(to_signed(-958,16));
ROM(2838) <= std_logic_vector(to_signed(-959,16));
ROM(2839) <= std_logic_vector(to_signed(-959,16));
ROM(2840) <= std_logic_vector(to_signed(-960,16));
ROM(2841) <= std_logic_vector(to_signed(-960,16));
ROM(2842) <= std_logic_vector(to_signed(-961,16));
ROM(2843) <= std_logic_vector(to_signed(-961,16));
ROM(2844) <= std_logic_vector(to_signed(-962,16));
ROM(2845) <= std_logic_vector(to_signed(-963,16));
ROM(2846) <= std_logic_vector(to_signed(-963,16));
ROM(2847) <= std_logic_vector(to_signed(-964,16));
ROM(2848) <= std_logic_vector(to_signed(-964,16));
ROM(2849) <= std_logic_vector(to_signed(-965,16));
ROM(2850) <= std_logic_vector(to_signed(-965,16));
ROM(2851) <= std_logic_vector(to_signed(-966,16));
ROM(2852) <= std_logic_vector(to_signed(-966,16));
ROM(2853) <= std_logic_vector(to_signed(-967,16));
ROM(2854) <= std_logic_vector(to_signed(-967,16));
ROM(2855) <= std_logic_vector(to_signed(-968,16));
ROM(2856) <= std_logic_vector(to_signed(-968,16));
ROM(2857) <= std_logic_vector(to_signed(-969,16));
ROM(2858) <= std_logic_vector(to_signed(-969,16));
ROM(2859) <= std_logic_vector(to_signed(-970,16));
ROM(2860) <= std_logic_vector(to_signed(-970,16));
ROM(2861) <= std_logic_vector(to_signed(-971,16));
ROM(2862) <= std_logic_vector(to_signed(-971,16));
ROM(2863) <= std_logic_vector(to_signed(-972,16));
ROM(2864) <= std_logic_vector(to_signed(-972,16));
ROM(2865) <= std_logic_vector(to_signed(-973,16));
ROM(2866) <= std_logic_vector(to_signed(-973,16));
ROM(2867) <= std_logic_vector(to_signed(-974,16));
ROM(2868) <= std_logic_vector(to_signed(-974,16));
ROM(2869) <= std_logic_vector(to_signed(-975,16));
ROM(2870) <= std_logic_vector(to_signed(-975,16));
ROM(2871) <= std_logic_vector(to_signed(-976,16));
ROM(2872) <= std_logic_vector(to_signed(-976,16));
ROM(2873) <= std_logic_vector(to_signed(-977,16));
ROM(2874) <= std_logic_vector(to_signed(-977,16));
ROM(2875) <= std_logic_vector(to_signed(-978,16));
ROM(2876) <= std_logic_vector(to_signed(-978,16));
ROM(2877) <= std_logic_vector(to_signed(-979,16));
ROM(2878) <= std_logic_vector(to_signed(-979,16));
ROM(2879) <= std_logic_vector(to_signed(-979,16));
ROM(2880) <= std_logic_vector(to_signed(-980,16));
ROM(2881) <= std_logic_vector(to_signed(-980,16));
ROM(2882) <= std_logic_vector(to_signed(-981,16));
ROM(2883) <= std_logic_vector(to_signed(-981,16));
ROM(2884) <= std_logic_vector(to_signed(-982,16));
ROM(2885) <= std_logic_vector(to_signed(-982,16));
ROM(2886) <= std_logic_vector(to_signed(-983,16));
ROM(2887) <= std_logic_vector(to_signed(-983,16));
ROM(2888) <= std_logic_vector(to_signed(-983,16));
ROM(2889) <= std_logic_vector(to_signed(-984,16));
ROM(2890) <= std_logic_vector(to_signed(-984,16));
ROM(2891) <= std_logic_vector(to_signed(-985,16));
ROM(2892) <= std_logic_vector(to_signed(-985,16));
ROM(2893) <= std_logic_vector(to_signed(-986,16));
ROM(2894) <= std_logic_vector(to_signed(-986,16));
ROM(2895) <= std_logic_vector(to_signed(-986,16));
ROM(2896) <= std_logic_vector(to_signed(-987,16));
ROM(2897) <= std_logic_vector(to_signed(-987,16));
ROM(2898) <= std_logic_vector(to_signed(-988,16));
ROM(2899) <= std_logic_vector(to_signed(-988,16));
ROM(2900) <= std_logic_vector(to_signed(-989,16));
ROM(2901) <= std_logic_vector(to_signed(-989,16));
ROM(2902) <= std_logic_vector(to_signed(-989,16));
ROM(2903) <= std_logic_vector(to_signed(-990,16));
ROM(2904) <= std_logic_vector(to_signed(-990,16));
ROM(2905) <= std_logic_vector(to_signed(-991,16));
ROM(2906) <= std_logic_vector(to_signed(-991,16));
ROM(2907) <= std_logic_vector(to_signed(-991,16));
ROM(2908) <= std_logic_vector(to_signed(-992,16));
ROM(2909) <= std_logic_vector(to_signed(-992,16));
ROM(2910) <= std_logic_vector(to_signed(-993,16));
ROM(2911) <= std_logic_vector(to_signed(-993,16));
ROM(2912) <= std_logic_vector(to_signed(-993,16));
ROM(2913) <= std_logic_vector(to_signed(-994,16));
ROM(2914) <= std_logic_vector(to_signed(-994,16));
ROM(2915) <= std_logic_vector(to_signed(-994,16));
ROM(2916) <= std_logic_vector(to_signed(-995,16));
ROM(2917) <= std_logic_vector(to_signed(-995,16));
ROM(2918) <= std_logic_vector(to_signed(-996,16));
ROM(2919) <= std_logic_vector(to_signed(-996,16));
ROM(2920) <= std_logic_vector(to_signed(-996,16));
ROM(2921) <= std_logic_vector(to_signed(-997,16));
ROM(2922) <= std_logic_vector(to_signed(-997,16));
ROM(2923) <= std_logic_vector(to_signed(-997,16));
ROM(2924) <= std_logic_vector(to_signed(-998,16));
ROM(2925) <= std_logic_vector(to_signed(-998,16));
ROM(2926) <= std_logic_vector(to_signed(-998,16));
ROM(2927) <= std_logic_vector(to_signed(-999,16));
ROM(2928) <= std_logic_vector(to_signed(-999,16));
ROM(2929) <= std_logic_vector(to_signed(-999,16));
ROM(2930) <= std_logic_vector(to_signed(-1000,16));
ROM(2931) <= std_logic_vector(to_signed(-1000,16));
ROM(2932) <= std_logic_vector(to_signed(-1000,16));
ROM(2933) <= std_logic_vector(to_signed(-1001,16));
ROM(2934) <= std_logic_vector(to_signed(-1001,16));
ROM(2935) <= std_logic_vector(to_signed(-1001,16));
ROM(2936) <= std_logic_vector(to_signed(-1002,16));
ROM(2937) <= std_logic_vector(to_signed(-1002,16));
ROM(2938) <= std_logic_vector(to_signed(-1002,16));
ROM(2939) <= std_logic_vector(to_signed(-1003,16));
ROM(2940) <= std_logic_vector(to_signed(-1003,16));
ROM(2941) <= std_logic_vector(to_signed(-1003,16));
ROM(2942) <= std_logic_vector(to_signed(-1004,16));
ROM(2943) <= std_logic_vector(to_signed(-1004,16));
ROM(2944) <= std_logic_vector(to_signed(-1004,16));
ROM(2945) <= std_logic_vector(to_signed(-1005,16));
ROM(2946) <= std_logic_vector(to_signed(-1005,16));
ROM(2947) <= std_logic_vector(to_signed(-1005,16));
ROM(2948) <= std_logic_vector(to_signed(-1006,16));
ROM(2949) <= std_logic_vector(to_signed(-1006,16));
ROM(2950) <= std_logic_vector(to_signed(-1006,16));
ROM(2951) <= std_logic_vector(to_signed(-1006,16));
ROM(2952) <= std_logic_vector(to_signed(-1007,16));
ROM(2953) <= std_logic_vector(to_signed(-1007,16));
ROM(2954) <= std_logic_vector(to_signed(-1007,16));
ROM(2955) <= std_logic_vector(to_signed(-1008,16));
ROM(2956) <= std_logic_vector(to_signed(-1008,16));
ROM(2957) <= std_logic_vector(to_signed(-1008,16));
ROM(2958) <= std_logic_vector(to_signed(-1008,16));
ROM(2959) <= std_logic_vector(to_signed(-1009,16));
ROM(2960) <= std_logic_vector(to_signed(-1009,16));
ROM(2961) <= std_logic_vector(to_signed(-1009,16));
ROM(2962) <= std_logic_vector(to_signed(-1009,16));
ROM(2963) <= std_logic_vector(to_signed(-1010,16));
ROM(2964) <= std_logic_vector(to_signed(-1010,16));
ROM(2965) <= std_logic_vector(to_signed(-1010,16));
ROM(2966) <= std_logic_vector(to_signed(-1010,16));
ROM(2967) <= std_logic_vector(to_signed(-1011,16));
ROM(2968) <= std_logic_vector(to_signed(-1011,16));
ROM(2969) <= std_logic_vector(to_signed(-1011,16));
ROM(2970) <= std_logic_vector(to_signed(-1011,16));
ROM(2971) <= std_logic_vector(to_signed(-1012,16));
ROM(2972) <= std_logic_vector(to_signed(-1012,16));
ROM(2973) <= std_logic_vector(to_signed(-1012,16));
ROM(2974) <= std_logic_vector(to_signed(-1012,16));
ROM(2975) <= std_logic_vector(to_signed(-1013,16));
ROM(2976) <= std_logic_vector(to_signed(-1013,16));
ROM(2977) <= std_logic_vector(to_signed(-1013,16));
ROM(2978) <= std_logic_vector(to_signed(-1013,16));
ROM(2979) <= std_logic_vector(to_signed(-1014,16));
ROM(2980) <= std_logic_vector(to_signed(-1014,16));
ROM(2981) <= std_logic_vector(to_signed(-1014,16));
ROM(2982) <= std_logic_vector(to_signed(-1014,16));
ROM(2983) <= std_logic_vector(to_signed(-1014,16));
ROM(2984) <= std_logic_vector(to_signed(-1015,16));
ROM(2985) <= std_logic_vector(to_signed(-1015,16));
ROM(2986) <= std_logic_vector(to_signed(-1015,16));
ROM(2987) <= std_logic_vector(to_signed(-1015,16));
ROM(2988) <= std_logic_vector(to_signed(-1016,16));
ROM(2989) <= std_logic_vector(to_signed(-1016,16));
ROM(2990) <= std_logic_vector(to_signed(-1016,16));
ROM(2991) <= std_logic_vector(to_signed(-1016,16));
ROM(2992) <= std_logic_vector(to_signed(-1016,16));
ROM(2993) <= std_logic_vector(to_signed(-1016,16));
ROM(2994) <= std_logic_vector(to_signed(-1017,16));
ROM(2995) <= std_logic_vector(to_signed(-1017,16));
ROM(2996) <= std_logic_vector(to_signed(-1017,16));
ROM(2997) <= std_logic_vector(to_signed(-1017,16));
ROM(2998) <= std_logic_vector(to_signed(-1017,16));
ROM(2999) <= std_logic_vector(to_signed(-1018,16));
ROM(3000) <= std_logic_vector(to_signed(-1018,16));
ROM(3001) <= std_logic_vector(to_signed(-1018,16));
ROM(3002) <= std_logic_vector(to_signed(-1018,16));
ROM(3003) <= std_logic_vector(to_signed(-1018,16));
ROM(3004) <= std_logic_vector(to_signed(-1018,16));
ROM(3005) <= std_logic_vector(to_signed(-1019,16));
ROM(3006) <= std_logic_vector(to_signed(-1019,16));
ROM(3007) <= std_logic_vector(to_signed(-1019,16));
ROM(3008) <= std_logic_vector(to_signed(-1019,16));
ROM(3009) <= std_logic_vector(to_signed(-1019,16));
ROM(3010) <= std_logic_vector(to_signed(-1019,16));
ROM(3011) <= std_logic_vector(to_signed(-1020,16));
ROM(3012) <= std_logic_vector(to_signed(-1020,16));
ROM(3013) <= std_logic_vector(to_signed(-1020,16));
ROM(3014) <= std_logic_vector(to_signed(-1020,16));
ROM(3015) <= std_logic_vector(to_signed(-1020,16));
ROM(3016) <= std_logic_vector(to_signed(-1020,16));
ROM(3017) <= std_logic_vector(to_signed(-1020,16));
ROM(3018) <= std_logic_vector(to_signed(-1020,16));
ROM(3019) <= std_logic_vector(to_signed(-1021,16));
ROM(3020) <= std_logic_vector(to_signed(-1021,16));
ROM(3021) <= std_logic_vector(to_signed(-1021,16));
ROM(3022) <= std_logic_vector(to_signed(-1021,16));
ROM(3023) <= std_logic_vector(to_signed(-1021,16));
ROM(3024) <= std_logic_vector(to_signed(-1021,16));
ROM(3025) <= std_logic_vector(to_signed(-1021,16));
ROM(3026) <= std_logic_vector(to_signed(-1021,16));
ROM(3027) <= std_logic_vector(to_signed(-1022,16));
ROM(3028) <= std_logic_vector(to_signed(-1022,16));
ROM(3029) <= std_logic_vector(to_signed(-1022,16));
ROM(3030) <= std_logic_vector(to_signed(-1022,16));
ROM(3031) <= std_logic_vector(to_signed(-1022,16));
ROM(3032) <= std_logic_vector(to_signed(-1022,16));
ROM(3033) <= std_logic_vector(to_signed(-1022,16));
ROM(3034) <= std_logic_vector(to_signed(-1022,16));
ROM(3035) <= std_logic_vector(to_signed(-1022,16));
ROM(3036) <= std_logic_vector(to_signed(-1022,16));
ROM(3037) <= std_logic_vector(to_signed(-1023,16));
ROM(3038) <= std_logic_vector(to_signed(-1023,16));
ROM(3039) <= std_logic_vector(to_signed(-1023,16));
ROM(3040) <= std_logic_vector(to_signed(-1023,16));
ROM(3041) <= std_logic_vector(to_signed(-1023,16));
ROM(3042) <= std_logic_vector(to_signed(-1023,16));
ROM(3043) <= std_logic_vector(to_signed(-1023,16));
ROM(3044) <= std_logic_vector(to_signed(-1023,16));
ROM(3045) <= std_logic_vector(to_signed(-1023,16));
ROM(3046) <= std_logic_vector(to_signed(-1023,16));
ROM(3047) <= std_logic_vector(to_signed(-1023,16));
ROM(3048) <= std_logic_vector(to_signed(-1023,16));
ROM(3049) <= std_logic_vector(to_signed(-1023,16));
ROM(3050) <= std_logic_vector(to_signed(-1023,16));
ROM(3051) <= std_logic_vector(to_signed(-1023,16));
ROM(3052) <= std_logic_vector(to_signed(-1024,16));
ROM(3053) <= std_logic_vector(to_signed(-1024,16));
ROM(3054) <= std_logic_vector(to_signed(-1024,16));
ROM(3055) <= std_logic_vector(to_signed(-1024,16));
ROM(3056) <= std_logic_vector(to_signed(-1024,16));
ROM(3057) <= std_logic_vector(to_signed(-1024,16));
ROM(3058) <= std_logic_vector(to_signed(-1024,16));
ROM(3059) <= std_logic_vector(to_signed(-1024,16));
ROM(3060) <= std_logic_vector(to_signed(-1024,16));
ROM(3061) <= std_logic_vector(to_signed(-1024,16));
ROM(3062) <= std_logic_vector(to_signed(-1024,16));
ROM(3063) <= std_logic_vector(to_signed(-1024,16));
ROM(3064) <= std_logic_vector(to_signed(-1024,16));
ROM(3065) <= std_logic_vector(to_signed(-1024,16));
ROM(3066) <= std_logic_vector(to_signed(-1024,16));
ROM(3067) <= std_logic_vector(to_signed(-1024,16));
ROM(3068) <= std_logic_vector(to_signed(-1024,16));
ROM(3069) <= std_logic_vector(to_signed(-1024,16));
ROM(3070) <= std_logic_vector(to_signed(-1024,16));
ROM(3071) <= std_logic_vector(to_signed(-1024,16));
ROM(3072) <= std_logic_vector(to_signed(-1024,16));
ROM(3073) <= std_logic_vector(to_signed(-1024,16));
ROM(3074) <= std_logic_vector(to_signed(-1024,16));
ROM(3075) <= std_logic_vector(to_signed(-1024,16));
ROM(3076) <= std_logic_vector(to_signed(-1024,16));
ROM(3077) <= std_logic_vector(to_signed(-1024,16));
ROM(3078) <= std_logic_vector(to_signed(-1024,16));
ROM(3079) <= std_logic_vector(to_signed(-1024,16));
ROM(3080) <= std_logic_vector(to_signed(-1024,16));
ROM(3081) <= std_logic_vector(to_signed(-1024,16));
ROM(3082) <= std_logic_vector(to_signed(-1024,16));
ROM(3083) <= std_logic_vector(to_signed(-1024,16));
ROM(3084) <= std_logic_vector(to_signed(-1024,16));
ROM(3085) <= std_logic_vector(to_signed(-1024,16));
ROM(3086) <= std_logic_vector(to_signed(-1024,16));
ROM(3087) <= std_logic_vector(to_signed(-1024,16));
ROM(3088) <= std_logic_vector(to_signed(-1024,16));
ROM(3089) <= std_logic_vector(to_signed(-1024,16));
ROM(3090) <= std_logic_vector(to_signed(-1024,16));
ROM(3091) <= std_logic_vector(to_signed(-1024,16));
ROM(3092) <= std_logic_vector(to_signed(-1024,16));
ROM(3093) <= std_logic_vector(to_signed(-1023,16));
ROM(3094) <= std_logic_vector(to_signed(-1023,16));
ROM(3095) <= std_logic_vector(to_signed(-1023,16));
ROM(3096) <= std_logic_vector(to_signed(-1023,16));
ROM(3097) <= std_logic_vector(to_signed(-1023,16));
ROM(3098) <= std_logic_vector(to_signed(-1023,16));
ROM(3099) <= std_logic_vector(to_signed(-1023,16));
ROM(3100) <= std_logic_vector(to_signed(-1023,16));
ROM(3101) <= std_logic_vector(to_signed(-1023,16));
ROM(3102) <= std_logic_vector(to_signed(-1023,16));
ROM(3103) <= std_logic_vector(to_signed(-1023,16));
ROM(3104) <= std_logic_vector(to_signed(-1023,16));
ROM(3105) <= std_logic_vector(to_signed(-1023,16));
ROM(3106) <= std_logic_vector(to_signed(-1023,16));
ROM(3107) <= std_logic_vector(to_signed(-1023,16));
ROM(3108) <= std_logic_vector(to_signed(-1022,16));
ROM(3109) <= std_logic_vector(to_signed(-1022,16));
ROM(3110) <= std_logic_vector(to_signed(-1022,16));
ROM(3111) <= std_logic_vector(to_signed(-1022,16));
ROM(3112) <= std_logic_vector(to_signed(-1022,16));
ROM(3113) <= std_logic_vector(to_signed(-1022,16));
ROM(3114) <= std_logic_vector(to_signed(-1022,16));
ROM(3115) <= std_logic_vector(to_signed(-1022,16));
ROM(3116) <= std_logic_vector(to_signed(-1022,16));
ROM(3117) <= std_logic_vector(to_signed(-1022,16));
ROM(3118) <= std_logic_vector(to_signed(-1021,16));
ROM(3119) <= std_logic_vector(to_signed(-1021,16));
ROM(3120) <= std_logic_vector(to_signed(-1021,16));
ROM(3121) <= std_logic_vector(to_signed(-1021,16));
ROM(3122) <= std_logic_vector(to_signed(-1021,16));
ROM(3123) <= std_logic_vector(to_signed(-1021,16));
ROM(3124) <= std_logic_vector(to_signed(-1021,16));
ROM(3125) <= std_logic_vector(to_signed(-1021,16));
ROM(3126) <= std_logic_vector(to_signed(-1020,16));
ROM(3127) <= std_logic_vector(to_signed(-1020,16));
ROM(3128) <= std_logic_vector(to_signed(-1020,16));
ROM(3129) <= std_logic_vector(to_signed(-1020,16));
ROM(3130) <= std_logic_vector(to_signed(-1020,16));
ROM(3131) <= std_logic_vector(to_signed(-1020,16));
ROM(3132) <= std_logic_vector(to_signed(-1020,16));
ROM(3133) <= std_logic_vector(to_signed(-1020,16));
ROM(3134) <= std_logic_vector(to_signed(-1019,16));
ROM(3135) <= std_logic_vector(to_signed(-1019,16));
ROM(3136) <= std_logic_vector(to_signed(-1019,16));
ROM(3137) <= std_logic_vector(to_signed(-1019,16));
ROM(3138) <= std_logic_vector(to_signed(-1019,16));
ROM(3139) <= std_logic_vector(to_signed(-1019,16));
ROM(3140) <= std_logic_vector(to_signed(-1018,16));
ROM(3141) <= std_logic_vector(to_signed(-1018,16));
ROM(3142) <= std_logic_vector(to_signed(-1018,16));
ROM(3143) <= std_logic_vector(to_signed(-1018,16));
ROM(3144) <= std_logic_vector(to_signed(-1018,16));
ROM(3145) <= std_logic_vector(to_signed(-1018,16));
ROM(3146) <= std_logic_vector(to_signed(-1017,16));
ROM(3147) <= std_logic_vector(to_signed(-1017,16));
ROM(3148) <= std_logic_vector(to_signed(-1017,16));
ROM(3149) <= std_logic_vector(to_signed(-1017,16));
ROM(3150) <= std_logic_vector(to_signed(-1017,16));
ROM(3151) <= std_logic_vector(to_signed(-1016,16));
ROM(3152) <= std_logic_vector(to_signed(-1016,16));
ROM(3153) <= std_logic_vector(to_signed(-1016,16));
ROM(3154) <= std_logic_vector(to_signed(-1016,16));
ROM(3155) <= std_logic_vector(to_signed(-1016,16));
ROM(3156) <= std_logic_vector(to_signed(-1016,16));
ROM(3157) <= std_logic_vector(to_signed(-1015,16));
ROM(3158) <= std_logic_vector(to_signed(-1015,16));
ROM(3159) <= std_logic_vector(to_signed(-1015,16));
ROM(3160) <= std_logic_vector(to_signed(-1015,16));
ROM(3161) <= std_logic_vector(to_signed(-1014,16));
ROM(3162) <= std_logic_vector(to_signed(-1014,16));
ROM(3163) <= std_logic_vector(to_signed(-1014,16));
ROM(3164) <= std_logic_vector(to_signed(-1014,16));
ROM(3165) <= std_logic_vector(to_signed(-1014,16));
ROM(3166) <= std_logic_vector(to_signed(-1013,16));
ROM(3167) <= std_logic_vector(to_signed(-1013,16));
ROM(3168) <= std_logic_vector(to_signed(-1013,16));
ROM(3169) <= std_logic_vector(to_signed(-1013,16));
ROM(3170) <= std_logic_vector(to_signed(-1012,16));
ROM(3171) <= std_logic_vector(to_signed(-1012,16));
ROM(3172) <= std_logic_vector(to_signed(-1012,16));
ROM(3173) <= std_logic_vector(to_signed(-1012,16));
ROM(3174) <= std_logic_vector(to_signed(-1011,16));
ROM(3175) <= std_logic_vector(to_signed(-1011,16));
ROM(3176) <= std_logic_vector(to_signed(-1011,16));
ROM(3177) <= std_logic_vector(to_signed(-1011,16));
ROM(3178) <= std_logic_vector(to_signed(-1010,16));
ROM(3179) <= std_logic_vector(to_signed(-1010,16));
ROM(3180) <= std_logic_vector(to_signed(-1010,16));
ROM(3181) <= std_logic_vector(to_signed(-1010,16));
ROM(3182) <= std_logic_vector(to_signed(-1009,16));
ROM(3183) <= std_logic_vector(to_signed(-1009,16));
ROM(3184) <= std_logic_vector(to_signed(-1009,16));
ROM(3185) <= std_logic_vector(to_signed(-1009,16));
ROM(3186) <= std_logic_vector(to_signed(-1008,16));
ROM(3187) <= std_logic_vector(to_signed(-1008,16));
ROM(3188) <= std_logic_vector(to_signed(-1008,16));
ROM(3189) <= std_logic_vector(to_signed(-1008,16));
ROM(3190) <= std_logic_vector(to_signed(-1007,16));
ROM(3191) <= std_logic_vector(to_signed(-1007,16));
ROM(3192) <= std_logic_vector(to_signed(-1007,16));
ROM(3193) <= std_logic_vector(to_signed(-1006,16));
ROM(3194) <= std_logic_vector(to_signed(-1006,16));
ROM(3195) <= std_logic_vector(to_signed(-1006,16));
ROM(3196) <= std_logic_vector(to_signed(-1006,16));
ROM(3197) <= std_logic_vector(to_signed(-1005,16));
ROM(3198) <= std_logic_vector(to_signed(-1005,16));
ROM(3199) <= std_logic_vector(to_signed(-1005,16));
ROM(3200) <= std_logic_vector(to_signed(-1004,16));
ROM(3201) <= std_logic_vector(to_signed(-1004,16));
ROM(3202) <= std_logic_vector(to_signed(-1004,16));
ROM(3203) <= std_logic_vector(to_signed(-1003,16));
ROM(3204) <= std_logic_vector(to_signed(-1003,16));
ROM(3205) <= std_logic_vector(to_signed(-1003,16));
ROM(3206) <= std_logic_vector(to_signed(-1002,16));
ROM(3207) <= std_logic_vector(to_signed(-1002,16));
ROM(3208) <= std_logic_vector(to_signed(-1002,16));
ROM(3209) <= std_logic_vector(to_signed(-1001,16));
ROM(3210) <= std_logic_vector(to_signed(-1001,16));
ROM(3211) <= std_logic_vector(to_signed(-1001,16));
ROM(3212) <= std_logic_vector(to_signed(-1000,16));
ROM(3213) <= std_logic_vector(to_signed(-1000,16));
ROM(3214) <= std_logic_vector(to_signed(-1000,16));
ROM(3215) <= std_logic_vector(to_signed(-999,16));
ROM(3216) <= std_logic_vector(to_signed(-999,16));
ROM(3217) <= std_logic_vector(to_signed(-999,16));
ROM(3218) <= std_logic_vector(to_signed(-998,16));
ROM(3219) <= std_logic_vector(to_signed(-998,16));
ROM(3220) <= std_logic_vector(to_signed(-998,16));
ROM(3221) <= std_logic_vector(to_signed(-997,16));
ROM(3222) <= std_logic_vector(to_signed(-997,16));
ROM(3223) <= std_logic_vector(to_signed(-997,16));
ROM(3224) <= std_logic_vector(to_signed(-996,16));
ROM(3225) <= std_logic_vector(to_signed(-996,16));
ROM(3226) <= std_logic_vector(to_signed(-996,16));
ROM(3227) <= std_logic_vector(to_signed(-995,16));
ROM(3228) <= std_logic_vector(to_signed(-995,16));
ROM(3229) <= std_logic_vector(to_signed(-994,16));
ROM(3230) <= std_logic_vector(to_signed(-994,16));
ROM(3231) <= std_logic_vector(to_signed(-994,16));
ROM(3232) <= std_logic_vector(to_signed(-993,16));
ROM(3233) <= std_logic_vector(to_signed(-993,16));
ROM(3234) <= std_logic_vector(to_signed(-993,16));
ROM(3235) <= std_logic_vector(to_signed(-992,16));
ROM(3236) <= std_logic_vector(to_signed(-992,16));
ROM(3237) <= std_logic_vector(to_signed(-991,16));
ROM(3238) <= std_logic_vector(to_signed(-991,16));
ROM(3239) <= std_logic_vector(to_signed(-991,16));
ROM(3240) <= std_logic_vector(to_signed(-990,16));
ROM(3241) <= std_logic_vector(to_signed(-990,16));
ROM(3242) <= std_logic_vector(to_signed(-989,16));
ROM(3243) <= std_logic_vector(to_signed(-989,16));
ROM(3244) <= std_logic_vector(to_signed(-989,16));
ROM(3245) <= std_logic_vector(to_signed(-988,16));
ROM(3246) <= std_logic_vector(to_signed(-988,16));
ROM(3247) <= std_logic_vector(to_signed(-987,16));
ROM(3248) <= std_logic_vector(to_signed(-987,16));
ROM(3249) <= std_logic_vector(to_signed(-986,16));
ROM(3250) <= std_logic_vector(to_signed(-986,16));
ROM(3251) <= std_logic_vector(to_signed(-986,16));
ROM(3252) <= std_logic_vector(to_signed(-985,16));
ROM(3253) <= std_logic_vector(to_signed(-985,16));
ROM(3254) <= std_logic_vector(to_signed(-984,16));
ROM(3255) <= std_logic_vector(to_signed(-984,16));
ROM(3256) <= std_logic_vector(to_signed(-983,16));
ROM(3257) <= std_logic_vector(to_signed(-983,16));
ROM(3258) <= std_logic_vector(to_signed(-983,16));
ROM(3259) <= std_logic_vector(to_signed(-982,16));
ROM(3260) <= std_logic_vector(to_signed(-982,16));
ROM(3261) <= std_logic_vector(to_signed(-981,16));
ROM(3262) <= std_logic_vector(to_signed(-981,16));
ROM(3263) <= std_logic_vector(to_signed(-980,16));
ROM(3264) <= std_logic_vector(to_signed(-980,16));
ROM(3265) <= std_logic_vector(to_signed(-979,16));
ROM(3266) <= std_logic_vector(to_signed(-979,16));
ROM(3267) <= std_logic_vector(to_signed(-979,16));
ROM(3268) <= std_logic_vector(to_signed(-978,16));
ROM(3269) <= std_logic_vector(to_signed(-978,16));
ROM(3270) <= std_logic_vector(to_signed(-977,16));
ROM(3271) <= std_logic_vector(to_signed(-977,16));
ROM(3272) <= std_logic_vector(to_signed(-976,16));
ROM(3273) <= std_logic_vector(to_signed(-976,16));
ROM(3274) <= std_logic_vector(to_signed(-975,16));
ROM(3275) <= std_logic_vector(to_signed(-975,16));
ROM(3276) <= std_logic_vector(to_signed(-974,16));
ROM(3277) <= std_logic_vector(to_signed(-974,16));
ROM(3278) <= std_logic_vector(to_signed(-973,16));
ROM(3279) <= std_logic_vector(to_signed(-973,16));
ROM(3280) <= std_logic_vector(to_signed(-972,16));
ROM(3281) <= std_logic_vector(to_signed(-972,16));
ROM(3282) <= std_logic_vector(to_signed(-971,16));
ROM(3283) <= std_logic_vector(to_signed(-971,16));
ROM(3284) <= std_logic_vector(to_signed(-970,16));
ROM(3285) <= std_logic_vector(to_signed(-970,16));
ROM(3286) <= std_logic_vector(to_signed(-969,16));
ROM(3287) <= std_logic_vector(to_signed(-969,16));
ROM(3288) <= std_logic_vector(to_signed(-968,16));
ROM(3289) <= std_logic_vector(to_signed(-968,16));
ROM(3290) <= std_logic_vector(to_signed(-967,16));
ROM(3291) <= std_logic_vector(to_signed(-967,16));
ROM(3292) <= std_logic_vector(to_signed(-966,16));
ROM(3293) <= std_logic_vector(to_signed(-966,16));
ROM(3294) <= std_logic_vector(to_signed(-965,16));
ROM(3295) <= std_logic_vector(to_signed(-965,16));
ROM(3296) <= std_logic_vector(to_signed(-964,16));
ROM(3297) <= std_logic_vector(to_signed(-964,16));
ROM(3298) <= std_logic_vector(to_signed(-963,16));
ROM(3299) <= std_logic_vector(to_signed(-963,16));
ROM(3300) <= std_logic_vector(to_signed(-962,16));
ROM(3301) <= std_logic_vector(to_signed(-961,16));
ROM(3302) <= std_logic_vector(to_signed(-961,16));
ROM(3303) <= std_logic_vector(to_signed(-960,16));
ROM(3304) <= std_logic_vector(to_signed(-960,16));
ROM(3305) <= std_logic_vector(to_signed(-959,16));
ROM(3306) <= std_logic_vector(to_signed(-959,16));
ROM(3307) <= std_logic_vector(to_signed(-958,16));
ROM(3308) <= std_logic_vector(to_signed(-958,16));
ROM(3309) <= std_logic_vector(to_signed(-957,16));
ROM(3310) <= std_logic_vector(to_signed(-957,16));
ROM(3311) <= std_logic_vector(to_signed(-956,16));
ROM(3312) <= std_logic_vector(to_signed(-955,16));
ROM(3313) <= std_logic_vector(to_signed(-955,16));
ROM(3314) <= std_logic_vector(to_signed(-954,16));
ROM(3315) <= std_logic_vector(to_signed(-954,16));
ROM(3316) <= std_logic_vector(to_signed(-953,16));
ROM(3317) <= std_logic_vector(to_signed(-953,16));
ROM(3318) <= std_logic_vector(to_signed(-952,16));
ROM(3319) <= std_logic_vector(to_signed(-951,16));
ROM(3320) <= std_logic_vector(to_signed(-951,16));
ROM(3321) <= std_logic_vector(to_signed(-950,16));
ROM(3322) <= std_logic_vector(to_signed(-950,16));
ROM(3323) <= std_logic_vector(to_signed(-949,16));
ROM(3324) <= std_logic_vector(to_signed(-948,16));
ROM(3325) <= std_logic_vector(to_signed(-948,16));
ROM(3326) <= std_logic_vector(to_signed(-947,16));
ROM(3327) <= std_logic_vector(to_signed(-947,16));
ROM(3328) <= std_logic_vector(to_signed(-946,16));
ROM(3329) <= std_logic_vector(to_signed(-945,16));
ROM(3330) <= std_logic_vector(to_signed(-945,16));
ROM(3331) <= std_logic_vector(to_signed(-944,16));
ROM(3332) <= std_logic_vector(to_signed(-944,16));
ROM(3333) <= std_logic_vector(to_signed(-943,16));
ROM(3334) <= std_logic_vector(to_signed(-942,16));
ROM(3335) <= std_logic_vector(to_signed(-942,16));
ROM(3336) <= std_logic_vector(to_signed(-941,16));
ROM(3337) <= std_logic_vector(to_signed(-941,16));
ROM(3338) <= std_logic_vector(to_signed(-940,16));
ROM(3339) <= std_logic_vector(to_signed(-939,16));
ROM(3340) <= std_logic_vector(to_signed(-939,16));
ROM(3341) <= std_logic_vector(to_signed(-938,16));
ROM(3342) <= std_logic_vector(to_signed(-937,16));
ROM(3343) <= std_logic_vector(to_signed(-937,16));
ROM(3344) <= std_logic_vector(to_signed(-936,16));
ROM(3345) <= std_logic_vector(to_signed(-936,16));
ROM(3346) <= std_logic_vector(to_signed(-935,16));
ROM(3347) <= std_logic_vector(to_signed(-934,16));
ROM(3348) <= std_logic_vector(to_signed(-934,16));
ROM(3349) <= std_logic_vector(to_signed(-933,16));
ROM(3350) <= std_logic_vector(to_signed(-932,16));
ROM(3351) <= std_logic_vector(to_signed(-932,16));
ROM(3352) <= std_logic_vector(to_signed(-931,16));
ROM(3353) <= std_logic_vector(to_signed(-930,16));
ROM(3354) <= std_logic_vector(to_signed(-930,16));
ROM(3355) <= std_logic_vector(to_signed(-929,16));
ROM(3356) <= std_logic_vector(to_signed(-928,16));
ROM(3357) <= std_logic_vector(to_signed(-928,16));
ROM(3358) <= std_logic_vector(to_signed(-927,16));
ROM(3359) <= std_logic_vector(to_signed(-926,16));
ROM(3360) <= std_logic_vector(to_signed(-926,16));
ROM(3361) <= std_logic_vector(to_signed(-925,16));
ROM(3362) <= std_logic_vector(to_signed(-924,16));
ROM(3363) <= std_logic_vector(to_signed(-924,16));
ROM(3364) <= std_logic_vector(to_signed(-923,16));
ROM(3365) <= std_logic_vector(to_signed(-922,16));
ROM(3366) <= std_logic_vector(to_signed(-922,16));
ROM(3367) <= std_logic_vector(to_signed(-921,16));
ROM(3368) <= std_logic_vector(to_signed(-920,16));
ROM(3369) <= std_logic_vector(to_signed(-920,16));
ROM(3370) <= std_logic_vector(to_signed(-919,16));
ROM(3371) <= std_logic_vector(to_signed(-918,16));
ROM(3372) <= std_logic_vector(to_signed(-917,16));
ROM(3373) <= std_logic_vector(to_signed(-917,16));
ROM(3374) <= std_logic_vector(to_signed(-916,16));
ROM(3375) <= std_logic_vector(to_signed(-915,16));
ROM(3376) <= std_logic_vector(to_signed(-915,16));
ROM(3377) <= std_logic_vector(to_signed(-914,16));
ROM(3378) <= std_logic_vector(to_signed(-913,16));
ROM(3379) <= std_logic_vector(to_signed(-913,16));
ROM(3380) <= std_logic_vector(to_signed(-912,16));
ROM(3381) <= std_logic_vector(to_signed(-911,16));
ROM(3382) <= std_logic_vector(to_signed(-910,16));
ROM(3383) <= std_logic_vector(to_signed(-910,16));
ROM(3384) <= std_logic_vector(to_signed(-909,16));
ROM(3385) <= std_logic_vector(to_signed(-908,16));
ROM(3386) <= std_logic_vector(to_signed(-907,16));
ROM(3387) <= std_logic_vector(to_signed(-907,16));
ROM(3388) <= std_logic_vector(to_signed(-906,16));
ROM(3389) <= std_logic_vector(to_signed(-905,16));
ROM(3390) <= std_logic_vector(to_signed(-905,16));
ROM(3391) <= std_logic_vector(to_signed(-904,16));
ROM(3392) <= std_logic_vector(to_signed(-903,16));
ROM(3393) <= std_logic_vector(to_signed(-902,16));
ROM(3394) <= std_logic_vector(to_signed(-902,16));
ROM(3395) <= std_logic_vector(to_signed(-901,16));
ROM(3396) <= std_logic_vector(to_signed(-900,16));
ROM(3397) <= std_logic_vector(to_signed(-899,16));
ROM(3398) <= std_logic_vector(to_signed(-899,16));
ROM(3399) <= std_logic_vector(to_signed(-898,16));
ROM(3400) <= std_logic_vector(to_signed(-897,16));
ROM(3401) <= std_logic_vector(to_signed(-896,16));
ROM(3402) <= std_logic_vector(to_signed(-896,16));
ROM(3403) <= std_logic_vector(to_signed(-895,16));
ROM(3404) <= std_logic_vector(to_signed(-894,16));
ROM(3405) <= std_logic_vector(to_signed(-893,16));
ROM(3406) <= std_logic_vector(to_signed(-893,16));
ROM(3407) <= std_logic_vector(to_signed(-892,16));
ROM(3408) <= std_logic_vector(to_signed(-891,16));
ROM(3409) <= std_logic_vector(to_signed(-890,16));
ROM(3410) <= std_logic_vector(to_signed(-889,16));
ROM(3411) <= std_logic_vector(to_signed(-889,16));
ROM(3412) <= std_logic_vector(to_signed(-888,16));
ROM(3413) <= std_logic_vector(to_signed(-887,16));
ROM(3414) <= std_logic_vector(to_signed(-886,16));
ROM(3415) <= std_logic_vector(to_signed(-885,16));
ROM(3416) <= std_logic_vector(to_signed(-885,16));
ROM(3417) <= std_logic_vector(to_signed(-884,16));
ROM(3418) <= std_logic_vector(to_signed(-883,16));
ROM(3419) <= std_logic_vector(to_signed(-882,16));
ROM(3420) <= std_logic_vector(to_signed(-882,16));
ROM(3421) <= std_logic_vector(to_signed(-881,16));
ROM(3422) <= std_logic_vector(to_signed(-880,16));
ROM(3423) <= std_logic_vector(to_signed(-879,16));
ROM(3424) <= std_logic_vector(to_signed(-878,16));
ROM(3425) <= std_logic_vector(to_signed(-878,16));
ROM(3426) <= std_logic_vector(to_signed(-877,16));
ROM(3427) <= std_logic_vector(to_signed(-876,16));
ROM(3428) <= std_logic_vector(to_signed(-875,16));
ROM(3429) <= std_logic_vector(to_signed(-874,16));
ROM(3430) <= std_logic_vector(to_signed(-873,16));
ROM(3431) <= std_logic_vector(to_signed(-873,16));
ROM(3432) <= std_logic_vector(to_signed(-872,16));
ROM(3433) <= std_logic_vector(to_signed(-871,16));
ROM(3434) <= std_logic_vector(to_signed(-870,16));
ROM(3435) <= std_logic_vector(to_signed(-869,16));
ROM(3436) <= std_logic_vector(to_signed(-868,16));
ROM(3437) <= std_logic_vector(to_signed(-868,16));
ROM(3438) <= std_logic_vector(to_signed(-867,16));
ROM(3439) <= std_logic_vector(to_signed(-866,16));
ROM(3440) <= std_logic_vector(to_signed(-865,16));
ROM(3441) <= std_logic_vector(to_signed(-864,16));
ROM(3442) <= std_logic_vector(to_signed(-863,16));
ROM(3443) <= std_logic_vector(to_signed(-863,16));
ROM(3444) <= std_logic_vector(to_signed(-862,16));
ROM(3445) <= std_logic_vector(to_signed(-861,16));
ROM(3446) <= std_logic_vector(to_signed(-860,16));
ROM(3447) <= std_logic_vector(to_signed(-859,16));
ROM(3448) <= std_logic_vector(to_signed(-858,16));
ROM(3449) <= std_logic_vector(to_signed(-857,16));
ROM(3450) <= std_logic_vector(to_signed(-857,16));
ROM(3451) <= std_logic_vector(to_signed(-856,16));
ROM(3452) <= std_logic_vector(to_signed(-855,16));
ROM(3453) <= std_logic_vector(to_signed(-854,16));
ROM(3454) <= std_logic_vector(to_signed(-853,16));
ROM(3455) <= std_logic_vector(to_signed(-852,16));
ROM(3456) <= std_logic_vector(to_signed(-851,16));
ROM(3457) <= std_logic_vector(to_signed(-851,16));
ROM(3458) <= std_logic_vector(to_signed(-850,16));
ROM(3459) <= std_logic_vector(to_signed(-849,16));
ROM(3460) <= std_logic_vector(to_signed(-848,16));
ROM(3461) <= std_logic_vector(to_signed(-847,16));
ROM(3462) <= std_logic_vector(to_signed(-846,16));
ROM(3463) <= std_logic_vector(to_signed(-845,16));
ROM(3464) <= std_logic_vector(to_signed(-844,16));
ROM(3465) <= std_logic_vector(to_signed(-843,16));
ROM(3466) <= std_logic_vector(to_signed(-843,16));
ROM(3467) <= std_logic_vector(to_signed(-842,16));
ROM(3468) <= std_logic_vector(to_signed(-841,16));
ROM(3469) <= std_logic_vector(to_signed(-840,16));
ROM(3470) <= std_logic_vector(to_signed(-839,16));
ROM(3471) <= std_logic_vector(to_signed(-838,16));
ROM(3472) <= std_logic_vector(to_signed(-837,16));
ROM(3473) <= std_logic_vector(to_signed(-836,16));
ROM(3474) <= std_logic_vector(to_signed(-835,16));
ROM(3475) <= std_logic_vector(to_signed(-834,16));
ROM(3476) <= std_logic_vector(to_signed(-834,16));
ROM(3477) <= std_logic_vector(to_signed(-833,16));
ROM(3478) <= std_logic_vector(to_signed(-832,16));
ROM(3479) <= std_logic_vector(to_signed(-831,16));
ROM(3480) <= std_logic_vector(to_signed(-830,16));
ROM(3481) <= std_logic_vector(to_signed(-829,16));
ROM(3482) <= std_logic_vector(to_signed(-828,16));
ROM(3483) <= std_logic_vector(to_signed(-827,16));
ROM(3484) <= std_logic_vector(to_signed(-826,16));
ROM(3485) <= std_logic_vector(to_signed(-825,16));
ROM(3486) <= std_logic_vector(to_signed(-824,16));
ROM(3487) <= std_logic_vector(to_signed(-823,16));
ROM(3488) <= std_logic_vector(to_signed(-822,16));
ROM(3489) <= std_logic_vector(to_signed(-822,16));
ROM(3490) <= std_logic_vector(to_signed(-821,16));
ROM(3491) <= std_logic_vector(to_signed(-820,16));
ROM(3492) <= std_logic_vector(to_signed(-819,16));
ROM(3493) <= std_logic_vector(to_signed(-818,16));
ROM(3494) <= std_logic_vector(to_signed(-817,16));
ROM(3495) <= std_logic_vector(to_signed(-816,16));
ROM(3496) <= std_logic_vector(to_signed(-815,16));
ROM(3497) <= std_logic_vector(to_signed(-814,16));
ROM(3498) <= std_logic_vector(to_signed(-813,16));
ROM(3499) <= std_logic_vector(to_signed(-812,16));
ROM(3500) <= std_logic_vector(to_signed(-811,16));
ROM(3501) <= std_logic_vector(to_signed(-810,16));
ROM(3502) <= std_logic_vector(to_signed(-809,16));
ROM(3503) <= std_logic_vector(to_signed(-808,16));
ROM(3504) <= std_logic_vector(to_signed(-807,16));
ROM(3505) <= std_logic_vector(to_signed(-806,16));
ROM(3506) <= std_logic_vector(to_signed(-805,16));
ROM(3507) <= std_logic_vector(to_signed(-804,16));
ROM(3508) <= std_logic_vector(to_signed(-803,16));
ROM(3509) <= std_logic_vector(to_signed(-802,16));
ROM(3510) <= std_logic_vector(to_signed(-801,16));
ROM(3511) <= std_logic_vector(to_signed(-800,16));
ROM(3512) <= std_logic_vector(to_signed(-799,16));
ROM(3513) <= std_logic_vector(to_signed(-798,16));
ROM(3514) <= std_logic_vector(to_signed(-798,16));
ROM(3515) <= std_logic_vector(to_signed(-797,16));
ROM(3516) <= std_logic_vector(to_signed(-796,16));
ROM(3517) <= std_logic_vector(to_signed(-795,16));
ROM(3518) <= std_logic_vector(to_signed(-794,16));
ROM(3519) <= std_logic_vector(to_signed(-793,16));
ROM(3520) <= std_logic_vector(to_signed(-792,16));
ROM(3521) <= std_logic_vector(to_signed(-791,16));
ROM(3522) <= std_logic_vector(to_signed(-790,16));
ROM(3523) <= std_logic_vector(to_signed(-789,16));
ROM(3524) <= std_logic_vector(to_signed(-788,16));
ROM(3525) <= std_logic_vector(to_signed(-787,16));
ROM(3526) <= std_logic_vector(to_signed(-786,16));
ROM(3527) <= std_logic_vector(to_signed(-785,16));
ROM(3528) <= std_logic_vector(to_signed(-784,16));
ROM(3529) <= std_logic_vector(to_signed(-783,16));
ROM(3530) <= std_logic_vector(to_signed(-782,16));
ROM(3531) <= std_logic_vector(to_signed(-780,16));
ROM(3532) <= std_logic_vector(to_signed(-779,16));
ROM(3533) <= std_logic_vector(to_signed(-778,16));
ROM(3534) <= std_logic_vector(to_signed(-777,16));
ROM(3535) <= std_logic_vector(to_signed(-776,16));
ROM(3536) <= std_logic_vector(to_signed(-775,16));
ROM(3537) <= std_logic_vector(to_signed(-774,16));
ROM(3538) <= std_logic_vector(to_signed(-773,16));
ROM(3539) <= std_logic_vector(to_signed(-772,16));
ROM(3540) <= std_logic_vector(to_signed(-771,16));
ROM(3541) <= std_logic_vector(to_signed(-770,16));
ROM(3542) <= std_logic_vector(to_signed(-769,16));
ROM(3543) <= std_logic_vector(to_signed(-768,16));
ROM(3544) <= std_logic_vector(to_signed(-767,16));
ROM(3545) <= std_logic_vector(to_signed(-766,16));
ROM(3546) <= std_logic_vector(to_signed(-765,16));
ROM(3547) <= std_logic_vector(to_signed(-764,16));
ROM(3548) <= std_logic_vector(to_signed(-763,16));
ROM(3549) <= std_logic_vector(to_signed(-762,16));
ROM(3550) <= std_logic_vector(to_signed(-761,16));
ROM(3551) <= std_logic_vector(to_signed(-760,16));
ROM(3552) <= std_logic_vector(to_signed(-759,16));
ROM(3553) <= std_logic_vector(to_signed(-758,16));
ROM(3554) <= std_logic_vector(to_signed(-757,16));
ROM(3555) <= std_logic_vector(to_signed(-756,16));
ROM(3556) <= std_logic_vector(to_signed(-755,16));
ROM(3557) <= std_logic_vector(to_signed(-753,16));
ROM(3558) <= std_logic_vector(to_signed(-752,16));
ROM(3559) <= std_logic_vector(to_signed(-751,16));
ROM(3560) <= std_logic_vector(to_signed(-750,16));
ROM(3561) <= std_logic_vector(to_signed(-749,16));
ROM(3562) <= std_logic_vector(to_signed(-748,16));
ROM(3563) <= std_logic_vector(to_signed(-747,16));
ROM(3564) <= std_logic_vector(to_signed(-746,16));
ROM(3565) <= std_logic_vector(to_signed(-745,16));
ROM(3566) <= std_logic_vector(to_signed(-744,16));
ROM(3567) <= std_logic_vector(to_signed(-743,16));
ROM(3568) <= std_logic_vector(to_signed(-742,16));
ROM(3569) <= std_logic_vector(to_signed(-741,16));
ROM(3570) <= std_logic_vector(to_signed(-739,16));
ROM(3571) <= std_logic_vector(to_signed(-738,16));
ROM(3572) <= std_logic_vector(to_signed(-737,16));
ROM(3573) <= std_logic_vector(to_signed(-736,16));
ROM(3574) <= std_logic_vector(to_signed(-735,16));
ROM(3575) <= std_logic_vector(to_signed(-734,16));
ROM(3576) <= std_logic_vector(to_signed(-733,16));
ROM(3577) <= std_logic_vector(to_signed(-732,16));
ROM(3578) <= std_logic_vector(to_signed(-731,16));
ROM(3579) <= std_logic_vector(to_signed(-730,16));
ROM(3580) <= std_logic_vector(to_signed(-729,16));
ROM(3581) <= std_logic_vector(to_signed(-727,16));
ROM(3582) <= std_logic_vector(to_signed(-726,16));
ROM(3583) <= std_logic_vector(to_signed(-725,16));
ROM(3584) <= std_logic_vector(to_signed(-724,16));
ROM(3585) <= std_logic_vector(to_signed(-723,16));
ROM(3586) <= std_logic_vector(to_signed(-722,16));
ROM(3587) <= std_logic_vector(to_signed(-721,16));
ROM(3588) <= std_logic_vector(to_signed(-720,16));
ROM(3589) <= std_logic_vector(to_signed(-719,16));
ROM(3590) <= std_logic_vector(to_signed(-717,16));
ROM(3591) <= std_logic_vector(to_signed(-716,16));
ROM(3592) <= std_logic_vector(to_signed(-715,16));
ROM(3593) <= std_logic_vector(to_signed(-714,16));
ROM(3594) <= std_logic_vector(to_signed(-713,16));
ROM(3595) <= std_logic_vector(to_signed(-712,16));
ROM(3596) <= std_logic_vector(to_signed(-711,16));
ROM(3597) <= std_logic_vector(to_signed(-709,16));
ROM(3598) <= std_logic_vector(to_signed(-708,16));
ROM(3599) <= std_logic_vector(to_signed(-707,16));
ROM(3600) <= std_logic_vector(to_signed(-706,16));
ROM(3601) <= std_logic_vector(to_signed(-705,16));
ROM(3602) <= std_logic_vector(to_signed(-704,16));
ROM(3603) <= std_logic_vector(to_signed(-703,16));
ROM(3604) <= std_logic_vector(to_signed(-702,16));
ROM(3605) <= std_logic_vector(to_signed(-700,16));
ROM(3606) <= std_logic_vector(to_signed(-699,16));
ROM(3607) <= std_logic_vector(to_signed(-698,16));
ROM(3608) <= std_logic_vector(to_signed(-697,16));
ROM(3609) <= std_logic_vector(to_signed(-696,16));
ROM(3610) <= std_logic_vector(to_signed(-695,16));
ROM(3611) <= std_logic_vector(to_signed(-693,16));
ROM(3612) <= std_logic_vector(to_signed(-692,16));
ROM(3613) <= std_logic_vector(to_signed(-691,16));
ROM(3614) <= std_logic_vector(to_signed(-690,16));
ROM(3615) <= std_logic_vector(to_signed(-689,16));
ROM(3616) <= std_logic_vector(to_signed(-688,16));
ROM(3617) <= std_logic_vector(to_signed(-687,16));
ROM(3618) <= std_logic_vector(to_signed(-685,16));
ROM(3619) <= std_logic_vector(to_signed(-684,16));
ROM(3620) <= std_logic_vector(to_signed(-683,16));
ROM(3621) <= std_logic_vector(to_signed(-682,16));
ROM(3622) <= std_logic_vector(to_signed(-681,16));
ROM(3623) <= std_logic_vector(to_signed(-679,16));
ROM(3624) <= std_logic_vector(to_signed(-678,16));
ROM(3625) <= std_logic_vector(to_signed(-677,16));
ROM(3626) <= std_logic_vector(to_signed(-676,16));
ROM(3627) <= std_logic_vector(to_signed(-675,16));
ROM(3628) <= std_logic_vector(to_signed(-674,16));
ROM(3629) <= std_logic_vector(to_signed(-672,16));
ROM(3630) <= std_logic_vector(to_signed(-671,16));
ROM(3631) <= std_logic_vector(to_signed(-670,16));
ROM(3632) <= std_logic_vector(to_signed(-669,16));
ROM(3633) <= std_logic_vector(to_signed(-668,16));
ROM(3634) <= std_logic_vector(to_signed(-666,16));
ROM(3635) <= std_logic_vector(to_signed(-665,16));
ROM(3636) <= std_logic_vector(to_signed(-664,16));
ROM(3637) <= std_logic_vector(to_signed(-663,16));
ROM(3638) <= std_logic_vector(to_signed(-662,16));
ROM(3639) <= std_logic_vector(to_signed(-660,16));
ROM(3640) <= std_logic_vector(to_signed(-659,16));
ROM(3641) <= std_logic_vector(to_signed(-658,16));
ROM(3642) <= std_logic_vector(to_signed(-657,16));
ROM(3643) <= std_logic_vector(to_signed(-656,16));
ROM(3644) <= std_logic_vector(to_signed(-654,16));
ROM(3645) <= std_logic_vector(to_signed(-653,16));
ROM(3646) <= std_logic_vector(to_signed(-652,16));
ROM(3647) <= std_logic_vector(to_signed(-651,16));
ROM(3648) <= std_logic_vector(to_signed(-650,16));
ROM(3649) <= std_logic_vector(to_signed(-648,16));
ROM(3650) <= std_logic_vector(to_signed(-647,16));
ROM(3651) <= std_logic_vector(to_signed(-646,16));
ROM(3652) <= std_logic_vector(to_signed(-645,16));
ROM(3653) <= std_logic_vector(to_signed(-644,16));
ROM(3654) <= std_logic_vector(to_signed(-642,16));
ROM(3655) <= std_logic_vector(to_signed(-641,16));
ROM(3656) <= std_logic_vector(to_signed(-640,16));
ROM(3657) <= std_logic_vector(to_signed(-639,16));
ROM(3658) <= std_logic_vector(to_signed(-637,16));
ROM(3659) <= std_logic_vector(to_signed(-636,16));
ROM(3660) <= std_logic_vector(to_signed(-635,16));
ROM(3661) <= std_logic_vector(to_signed(-634,16));
ROM(3662) <= std_logic_vector(to_signed(-632,16));
ROM(3663) <= std_logic_vector(to_signed(-631,16));
ROM(3664) <= std_logic_vector(to_signed(-630,16));
ROM(3665) <= std_logic_vector(to_signed(-629,16));
ROM(3666) <= std_logic_vector(to_signed(-628,16));
ROM(3667) <= std_logic_vector(to_signed(-626,16));
ROM(3668) <= std_logic_vector(to_signed(-625,16));
ROM(3669) <= std_logic_vector(to_signed(-624,16));
ROM(3670) <= std_logic_vector(to_signed(-623,16));
ROM(3671) <= std_logic_vector(to_signed(-621,16));
ROM(3672) <= std_logic_vector(to_signed(-620,16));
ROM(3673) <= std_logic_vector(to_signed(-619,16));
ROM(3674) <= std_logic_vector(to_signed(-618,16));
ROM(3675) <= std_logic_vector(to_signed(-616,16));
ROM(3676) <= std_logic_vector(to_signed(-615,16));
ROM(3677) <= std_logic_vector(to_signed(-614,16));
ROM(3678) <= std_logic_vector(to_signed(-613,16));
ROM(3679) <= std_logic_vector(to_signed(-611,16));
ROM(3680) <= std_logic_vector(to_signed(-610,16));
ROM(3681) <= std_logic_vector(to_signed(-609,16));
ROM(3682) <= std_logic_vector(to_signed(-607,16));
ROM(3683) <= std_logic_vector(to_signed(-606,16));
ROM(3684) <= std_logic_vector(to_signed(-605,16));
ROM(3685) <= std_logic_vector(to_signed(-604,16));
ROM(3686) <= std_logic_vector(to_signed(-602,16));
ROM(3687) <= std_logic_vector(to_signed(-601,16));
ROM(3688) <= std_logic_vector(to_signed(-600,16));
ROM(3689) <= std_logic_vector(to_signed(-599,16));
ROM(3690) <= std_logic_vector(to_signed(-597,16));
ROM(3691) <= std_logic_vector(to_signed(-596,16));
ROM(3692) <= std_logic_vector(to_signed(-595,16));
ROM(3693) <= std_logic_vector(to_signed(-593,16));
ROM(3694) <= std_logic_vector(to_signed(-592,16));
ROM(3695) <= std_logic_vector(to_signed(-591,16));
ROM(3696) <= std_logic_vector(to_signed(-590,16));
ROM(3697) <= std_logic_vector(to_signed(-588,16));
ROM(3698) <= std_logic_vector(to_signed(-587,16));
ROM(3699) <= std_logic_vector(to_signed(-586,16));
ROM(3700) <= std_logic_vector(to_signed(-584,16));
ROM(3701) <= std_logic_vector(to_signed(-583,16));
ROM(3702) <= std_logic_vector(to_signed(-582,16));
ROM(3703) <= std_logic_vector(to_signed(-581,16));
ROM(3704) <= std_logic_vector(to_signed(-579,16));
ROM(3705) <= std_logic_vector(to_signed(-578,16));
ROM(3706) <= std_logic_vector(to_signed(-577,16));
ROM(3707) <= std_logic_vector(to_signed(-575,16));
ROM(3708) <= std_logic_vector(to_signed(-574,16));
ROM(3709) <= std_logic_vector(to_signed(-573,16));
ROM(3710) <= std_logic_vector(to_signed(-572,16));
ROM(3711) <= std_logic_vector(to_signed(-570,16));
ROM(3712) <= std_logic_vector(to_signed(-569,16));
ROM(3713) <= std_logic_vector(to_signed(-568,16));
ROM(3714) <= std_logic_vector(to_signed(-566,16));
ROM(3715) <= std_logic_vector(to_signed(-565,16));
ROM(3716) <= std_logic_vector(to_signed(-564,16));
ROM(3717) <= std_logic_vector(to_signed(-562,16));
ROM(3718) <= std_logic_vector(to_signed(-561,16));
ROM(3719) <= std_logic_vector(to_signed(-560,16));
ROM(3720) <= std_logic_vector(to_signed(-558,16));
ROM(3721) <= std_logic_vector(to_signed(-557,16));
ROM(3722) <= std_logic_vector(to_signed(-556,16));
ROM(3723) <= std_logic_vector(to_signed(-554,16));
ROM(3724) <= std_logic_vector(to_signed(-553,16));
ROM(3725) <= std_logic_vector(to_signed(-552,16));
ROM(3726) <= std_logic_vector(to_signed(-550,16));
ROM(3727) <= std_logic_vector(to_signed(-549,16));
ROM(3728) <= std_logic_vector(to_signed(-548,16));
ROM(3729) <= std_logic_vector(to_signed(-547,16));
ROM(3730) <= std_logic_vector(to_signed(-545,16));
ROM(3731) <= std_logic_vector(to_signed(-544,16));
ROM(3732) <= std_logic_vector(to_signed(-543,16));
ROM(3733) <= std_logic_vector(to_signed(-541,16));
ROM(3734) <= std_logic_vector(to_signed(-540,16));
ROM(3735) <= std_logic_vector(to_signed(-539,16));
ROM(3736) <= std_logic_vector(to_signed(-537,16));
ROM(3737) <= std_logic_vector(to_signed(-536,16));
ROM(3738) <= std_logic_vector(to_signed(-535,16));
ROM(3739) <= std_logic_vector(to_signed(-533,16));
ROM(3740) <= std_logic_vector(to_signed(-532,16));
ROM(3741) <= std_logic_vector(to_signed(-530,16));
ROM(3742) <= std_logic_vector(to_signed(-529,16));
ROM(3743) <= std_logic_vector(to_signed(-528,16));
ROM(3744) <= std_logic_vector(to_signed(-526,16));
ROM(3745) <= std_logic_vector(to_signed(-525,16));
ROM(3746) <= std_logic_vector(to_signed(-524,16));
ROM(3747) <= std_logic_vector(to_signed(-522,16));
ROM(3748) <= std_logic_vector(to_signed(-521,16));
ROM(3749) <= std_logic_vector(to_signed(-520,16));
ROM(3750) <= std_logic_vector(to_signed(-518,16));
ROM(3751) <= std_logic_vector(to_signed(-517,16));
ROM(3752) <= std_logic_vector(to_signed(-516,16));
ROM(3753) <= std_logic_vector(to_signed(-514,16));
ROM(3754) <= std_logic_vector(to_signed(-513,16));
ROM(3755) <= std_logic_vector(to_signed(-512,16));
ROM(3756) <= std_logic_vector(to_signed(-510,16));
ROM(3757) <= std_logic_vector(to_signed(-509,16));
ROM(3758) <= std_logic_vector(to_signed(-507,16));
ROM(3759) <= std_logic_vector(to_signed(-506,16));
ROM(3760) <= std_logic_vector(to_signed(-505,16));
ROM(3761) <= std_logic_vector(to_signed(-503,16));
ROM(3762) <= std_logic_vector(to_signed(-502,16));
ROM(3763) <= std_logic_vector(to_signed(-501,16));
ROM(3764) <= std_logic_vector(to_signed(-499,16));
ROM(3765) <= std_logic_vector(to_signed(-498,16));
ROM(3766) <= std_logic_vector(to_signed(-497,16));
ROM(3767) <= std_logic_vector(to_signed(-495,16));
ROM(3768) <= std_logic_vector(to_signed(-494,16));
ROM(3769) <= std_logic_vector(to_signed(-492,16));
ROM(3770) <= std_logic_vector(to_signed(-491,16));
ROM(3771) <= std_logic_vector(to_signed(-490,16));
ROM(3772) <= std_logic_vector(to_signed(-488,16));
ROM(3773) <= std_logic_vector(to_signed(-487,16));
ROM(3774) <= std_logic_vector(to_signed(-485,16));
ROM(3775) <= std_logic_vector(to_signed(-484,16));
ROM(3776) <= std_logic_vector(to_signed(-483,16));
ROM(3777) <= std_logic_vector(to_signed(-481,16));
ROM(3778) <= std_logic_vector(to_signed(-480,16));
ROM(3779) <= std_logic_vector(to_signed(-479,16));
ROM(3780) <= std_logic_vector(to_signed(-477,16));
ROM(3781) <= std_logic_vector(to_signed(-476,16));
ROM(3782) <= std_logic_vector(to_signed(-474,16));
ROM(3783) <= std_logic_vector(to_signed(-473,16));
ROM(3784) <= std_logic_vector(to_signed(-472,16));
ROM(3785) <= std_logic_vector(to_signed(-470,16));
ROM(3786) <= std_logic_vector(to_signed(-469,16));
ROM(3787) <= std_logic_vector(to_signed(-467,16));
ROM(3788) <= std_logic_vector(to_signed(-466,16));
ROM(3789) <= std_logic_vector(to_signed(-465,16));
ROM(3790) <= std_logic_vector(to_signed(-463,16));
ROM(3791) <= std_logic_vector(to_signed(-462,16));
ROM(3792) <= std_logic_vector(to_signed(-460,16));
ROM(3793) <= std_logic_vector(to_signed(-459,16));
ROM(3794) <= std_logic_vector(to_signed(-458,16));
ROM(3795) <= std_logic_vector(to_signed(-456,16));
ROM(3796) <= std_logic_vector(to_signed(-455,16));
ROM(3797) <= std_logic_vector(to_signed(-453,16));
ROM(3798) <= std_logic_vector(to_signed(-452,16));
ROM(3799) <= std_logic_vector(to_signed(-451,16));
ROM(3800) <= std_logic_vector(to_signed(-449,16));
ROM(3801) <= std_logic_vector(to_signed(-448,16));
ROM(3802) <= std_logic_vector(to_signed(-446,16));
ROM(3803) <= std_logic_vector(to_signed(-445,16));
ROM(3804) <= std_logic_vector(to_signed(-443,16));
ROM(3805) <= std_logic_vector(to_signed(-442,16));
ROM(3806) <= std_logic_vector(to_signed(-441,16));
ROM(3807) <= std_logic_vector(to_signed(-439,16));
ROM(3808) <= std_logic_vector(to_signed(-438,16));
ROM(3809) <= std_logic_vector(to_signed(-436,16));
ROM(3810) <= std_logic_vector(to_signed(-435,16));
ROM(3811) <= std_logic_vector(to_signed(-434,16));
ROM(3812) <= std_logic_vector(to_signed(-432,16));
ROM(3813) <= std_logic_vector(to_signed(-431,16));
ROM(3814) <= std_logic_vector(to_signed(-429,16));
ROM(3815) <= std_logic_vector(to_signed(-428,16));
ROM(3816) <= std_logic_vector(to_signed(-426,16));
ROM(3817) <= std_logic_vector(to_signed(-425,16));
ROM(3818) <= std_logic_vector(to_signed(-424,16));
ROM(3819) <= std_logic_vector(to_signed(-422,16));
ROM(3820) <= std_logic_vector(to_signed(-421,16));
ROM(3821) <= std_logic_vector(to_signed(-419,16));
ROM(3822) <= std_logic_vector(to_signed(-418,16));
ROM(3823) <= std_logic_vector(to_signed(-416,16));
ROM(3824) <= std_logic_vector(to_signed(-415,16));
ROM(3825) <= std_logic_vector(to_signed(-414,16));
ROM(3826) <= std_logic_vector(to_signed(-412,16));
ROM(3827) <= std_logic_vector(to_signed(-411,16));
ROM(3828) <= std_logic_vector(to_signed(-409,16));
ROM(3829) <= std_logic_vector(to_signed(-408,16));
ROM(3830) <= std_logic_vector(to_signed(-406,16));
ROM(3831) <= std_logic_vector(to_signed(-405,16));
ROM(3832) <= std_logic_vector(to_signed(-403,16));
ROM(3833) <= std_logic_vector(to_signed(-402,16));
ROM(3834) <= std_logic_vector(to_signed(-401,16));
ROM(3835) <= std_logic_vector(to_signed(-399,16));
ROM(3836) <= std_logic_vector(to_signed(-398,16));
ROM(3837) <= std_logic_vector(to_signed(-396,16));
ROM(3838) <= std_logic_vector(to_signed(-395,16));
ROM(3839) <= std_logic_vector(to_signed(-393,16));
ROM(3840) <= std_logic_vector(to_signed(-392,16));
ROM(3841) <= std_logic_vector(to_signed(-390,16));
ROM(3842) <= std_logic_vector(to_signed(-389,16));
ROM(3843) <= std_logic_vector(to_signed(-388,16));
ROM(3844) <= std_logic_vector(to_signed(-386,16));
ROM(3845) <= std_logic_vector(to_signed(-385,16));
ROM(3846) <= std_logic_vector(to_signed(-383,16));
ROM(3847) <= std_logic_vector(to_signed(-382,16));
ROM(3848) <= std_logic_vector(to_signed(-380,16));
ROM(3849) <= std_logic_vector(to_signed(-379,16));
ROM(3850) <= std_logic_vector(to_signed(-377,16));
ROM(3851) <= std_logic_vector(to_signed(-376,16));
ROM(3852) <= std_logic_vector(to_signed(-374,16));
ROM(3853) <= std_logic_vector(to_signed(-373,16));
ROM(3854) <= std_logic_vector(to_signed(-371,16));
ROM(3855) <= std_logic_vector(to_signed(-370,16));
ROM(3856) <= std_logic_vector(to_signed(-369,16));
ROM(3857) <= std_logic_vector(to_signed(-367,16));
ROM(3858) <= std_logic_vector(to_signed(-366,16));
ROM(3859) <= std_logic_vector(to_signed(-364,16));
ROM(3860) <= std_logic_vector(to_signed(-363,16));
ROM(3861) <= std_logic_vector(to_signed(-361,16));
ROM(3862) <= std_logic_vector(to_signed(-360,16));
ROM(3863) <= std_logic_vector(to_signed(-358,16));
ROM(3864) <= std_logic_vector(to_signed(-357,16));
ROM(3865) <= std_logic_vector(to_signed(-355,16));
ROM(3866) <= std_logic_vector(to_signed(-354,16));
ROM(3867) <= std_logic_vector(to_signed(-352,16));
ROM(3868) <= std_logic_vector(to_signed(-351,16));
ROM(3869) <= std_logic_vector(to_signed(-349,16));
ROM(3870) <= std_logic_vector(to_signed(-348,16));
ROM(3871) <= std_logic_vector(to_signed(-346,16));
ROM(3872) <= std_logic_vector(to_signed(-345,16));
ROM(3873) <= std_logic_vector(to_signed(-343,16));
ROM(3874) <= std_logic_vector(to_signed(-342,16));
ROM(3875) <= std_logic_vector(to_signed(-341,16));
ROM(3876) <= std_logic_vector(to_signed(-339,16));
ROM(3877) <= std_logic_vector(to_signed(-338,16));
ROM(3878) <= std_logic_vector(to_signed(-336,16));
ROM(3879) <= std_logic_vector(to_signed(-335,16));
ROM(3880) <= std_logic_vector(to_signed(-333,16));
ROM(3881) <= std_logic_vector(to_signed(-332,16));
ROM(3882) <= std_logic_vector(to_signed(-330,16));
ROM(3883) <= std_logic_vector(to_signed(-329,16));
ROM(3884) <= std_logic_vector(to_signed(-327,16));
ROM(3885) <= std_logic_vector(to_signed(-326,16));
ROM(3886) <= std_logic_vector(to_signed(-324,16));
ROM(3887) <= std_logic_vector(to_signed(-323,16));
ROM(3888) <= std_logic_vector(to_signed(-321,16));
ROM(3889) <= std_logic_vector(to_signed(-320,16));
ROM(3890) <= std_logic_vector(to_signed(-318,16));
ROM(3891) <= std_logic_vector(to_signed(-317,16));
ROM(3892) <= std_logic_vector(to_signed(-315,16));
ROM(3893) <= std_logic_vector(to_signed(-314,16));
ROM(3894) <= std_logic_vector(to_signed(-312,16));
ROM(3895) <= std_logic_vector(to_signed(-311,16));
ROM(3896) <= std_logic_vector(to_signed(-309,16));
ROM(3897) <= std_logic_vector(to_signed(-308,16));
ROM(3898) <= std_logic_vector(to_signed(-306,16));
ROM(3899) <= std_logic_vector(to_signed(-305,16));
ROM(3900) <= std_logic_vector(to_signed(-303,16));
ROM(3901) <= std_logic_vector(to_signed(-302,16));
ROM(3902) <= std_logic_vector(to_signed(-300,16));
ROM(3903) <= std_logic_vector(to_signed(-299,16));
ROM(3904) <= std_logic_vector(to_signed(-297,16));
ROM(3905) <= std_logic_vector(to_signed(-296,16));
ROM(3906) <= std_logic_vector(to_signed(-294,16));
ROM(3907) <= std_logic_vector(to_signed(-293,16));
ROM(3908) <= std_logic_vector(to_signed(-291,16));
ROM(3909) <= std_logic_vector(to_signed(-290,16));
ROM(3910) <= std_logic_vector(to_signed(-288,16));
ROM(3911) <= std_logic_vector(to_signed(-287,16));
ROM(3912) <= std_logic_vector(to_signed(-285,16));
ROM(3913) <= std_logic_vector(to_signed(-284,16));
ROM(3914) <= std_logic_vector(to_signed(-282,16));
ROM(3915) <= std_logic_vector(to_signed(-281,16));
ROM(3916) <= std_logic_vector(to_signed(-279,16));
ROM(3917) <= std_logic_vector(to_signed(-278,16));
ROM(3918) <= std_logic_vector(to_signed(-276,16));
ROM(3919) <= std_logic_vector(to_signed(-275,16));
ROM(3920) <= std_logic_vector(to_signed(-273,16));
ROM(3921) <= std_logic_vector(to_signed(-272,16));
ROM(3922) <= std_logic_vector(to_signed(-270,16));
ROM(3923) <= std_logic_vector(to_signed(-269,16));
ROM(3924) <= std_logic_vector(to_signed(-267,16));
ROM(3925) <= std_logic_vector(to_signed(-266,16));
ROM(3926) <= std_logic_vector(to_signed(-264,16));
ROM(3927) <= std_logic_vector(to_signed(-263,16));
ROM(3928) <= std_logic_vector(to_signed(-261,16));
ROM(3929) <= std_logic_vector(to_signed(-259,16));
ROM(3930) <= std_logic_vector(to_signed(-258,16));
ROM(3931) <= std_logic_vector(to_signed(-256,16));
ROM(3932) <= std_logic_vector(to_signed(-255,16));
ROM(3933) <= std_logic_vector(to_signed(-253,16));
ROM(3934) <= std_logic_vector(to_signed(-252,16));
ROM(3935) <= std_logic_vector(to_signed(-250,16));
ROM(3936) <= std_logic_vector(to_signed(-249,16));
ROM(3937) <= std_logic_vector(to_signed(-247,16));
ROM(3938) <= std_logic_vector(to_signed(-246,16));
ROM(3939) <= std_logic_vector(to_signed(-244,16));
ROM(3940) <= std_logic_vector(to_signed(-243,16));
ROM(3941) <= std_logic_vector(to_signed(-241,16));
ROM(3942) <= std_logic_vector(to_signed(-240,16));
ROM(3943) <= std_logic_vector(to_signed(-238,16));
ROM(3944) <= std_logic_vector(to_signed(-237,16));
ROM(3945) <= std_logic_vector(to_signed(-235,16));
ROM(3946) <= std_logic_vector(to_signed(-234,16));
ROM(3947) <= std_logic_vector(to_signed(-232,16));
ROM(3948) <= std_logic_vector(to_signed(-230,16));
ROM(3949) <= std_logic_vector(to_signed(-229,16));
ROM(3950) <= std_logic_vector(to_signed(-227,16));
ROM(3951) <= std_logic_vector(to_signed(-226,16));
ROM(3952) <= std_logic_vector(to_signed(-224,16));
ROM(3953) <= std_logic_vector(to_signed(-223,16));
ROM(3954) <= std_logic_vector(to_signed(-221,16));
ROM(3955) <= std_logic_vector(to_signed(-220,16));
ROM(3956) <= std_logic_vector(to_signed(-218,16));
ROM(3957) <= std_logic_vector(to_signed(-217,16));
ROM(3958) <= std_logic_vector(to_signed(-215,16));
ROM(3959) <= std_logic_vector(to_signed(-214,16));
ROM(3960) <= std_logic_vector(to_signed(-212,16));
ROM(3961) <= std_logic_vector(to_signed(-211,16));
ROM(3962) <= std_logic_vector(to_signed(-209,16));
ROM(3963) <= std_logic_vector(to_signed(-207,16));
ROM(3964) <= std_logic_vector(to_signed(-206,16));
ROM(3965) <= std_logic_vector(to_signed(-204,16));
ROM(3966) <= std_logic_vector(to_signed(-203,16));
ROM(3967) <= std_logic_vector(to_signed(-201,16));
ROM(3968) <= std_logic_vector(to_signed(-200,16));
ROM(3969) <= std_logic_vector(to_signed(-198,16));
ROM(3970) <= std_logic_vector(to_signed(-197,16));
ROM(3971) <= std_logic_vector(to_signed(-195,16));
ROM(3972) <= std_logic_vector(to_signed(-194,16));
ROM(3973) <= std_logic_vector(to_signed(-192,16));
ROM(3974) <= std_logic_vector(to_signed(-191,16));
ROM(3975) <= std_logic_vector(to_signed(-189,16));
ROM(3976) <= std_logic_vector(to_signed(-187,16));
ROM(3977) <= std_logic_vector(to_signed(-186,16));
ROM(3978) <= std_logic_vector(to_signed(-184,16));
ROM(3979) <= std_logic_vector(to_signed(-183,16));
ROM(3980) <= std_logic_vector(to_signed(-181,16));
ROM(3981) <= std_logic_vector(to_signed(-180,16));
ROM(3982) <= std_logic_vector(to_signed(-178,16));
ROM(3983) <= std_logic_vector(to_signed(-177,16));
ROM(3984) <= std_logic_vector(to_signed(-175,16));
ROM(3985) <= std_logic_vector(to_signed(-174,16));
ROM(3986) <= std_logic_vector(to_signed(-172,16));
ROM(3987) <= std_logic_vector(to_signed(-170,16));
ROM(3988) <= std_logic_vector(to_signed(-169,16));
ROM(3989) <= std_logic_vector(to_signed(-167,16));
ROM(3990) <= std_logic_vector(to_signed(-166,16));
ROM(3991) <= std_logic_vector(to_signed(-164,16));
ROM(3992) <= std_logic_vector(to_signed(-163,16));
ROM(3993) <= std_logic_vector(to_signed(-161,16));
ROM(3994) <= std_logic_vector(to_signed(-160,16));
ROM(3995) <= std_logic_vector(to_signed(-158,16));
ROM(3996) <= std_logic_vector(to_signed(-156,16));
ROM(3997) <= std_logic_vector(to_signed(-155,16));
ROM(3998) <= std_logic_vector(to_signed(-153,16));
ROM(3999) <= std_logic_vector(to_signed(-152,16));
ROM(4000) <= std_logic_vector(to_signed(-150,16));
ROM(4001) <= std_logic_vector(to_signed(-149,16));
ROM(4002) <= std_logic_vector(to_signed(-147,16));
ROM(4003) <= std_logic_vector(to_signed(-146,16));
ROM(4004) <= std_logic_vector(to_signed(-144,16));
ROM(4005) <= std_logic_vector(to_signed(-142,16));
ROM(4006) <= std_logic_vector(to_signed(-141,16));
ROM(4007) <= std_logic_vector(to_signed(-139,16));
ROM(4008) <= std_logic_vector(to_signed(-138,16));
ROM(4009) <= std_logic_vector(to_signed(-136,16));
ROM(4010) <= std_logic_vector(to_signed(-135,16));
ROM(4011) <= std_logic_vector(to_signed(-133,16));
ROM(4012) <= std_logic_vector(to_signed(-132,16));
ROM(4013) <= std_logic_vector(to_signed(-130,16));
ROM(4014) <= std_logic_vector(to_signed(-128,16));
ROM(4015) <= std_logic_vector(to_signed(-127,16));
ROM(4016) <= std_logic_vector(to_signed(-125,16));
ROM(4017) <= std_logic_vector(to_signed(-124,16));
ROM(4018) <= std_logic_vector(to_signed(-122,16));
ROM(4019) <= std_logic_vector(to_signed(-121,16));
ROM(4020) <= std_logic_vector(to_signed(-119,16));
ROM(4021) <= std_logic_vector(to_signed(-118,16));
ROM(4022) <= std_logic_vector(to_signed(-116,16));
ROM(4023) <= std_logic_vector(to_signed(-114,16));
ROM(4024) <= std_logic_vector(to_signed(-113,16));
ROM(4025) <= std_logic_vector(to_signed(-111,16));
ROM(4026) <= std_logic_vector(to_signed(-110,16));
ROM(4027) <= std_logic_vector(to_signed(-108,16));
ROM(4028) <= std_logic_vector(to_signed(-107,16));
ROM(4029) <= std_logic_vector(to_signed(-105,16));
ROM(4030) <= std_logic_vector(to_signed(-103,16));
ROM(4031) <= std_logic_vector(to_signed(-102,16));
ROM(4032) <= std_logic_vector(to_signed(-100,16));
ROM(4033) <= std_logic_vector(to_signed(-99,16));
ROM(4034) <= std_logic_vector(to_signed(-97,16));
ROM(4035) <= std_logic_vector(to_signed(-96,16));
ROM(4036) <= std_logic_vector(to_signed(-94,16));
ROM(4037) <= std_logic_vector(to_signed(-93,16));
ROM(4038) <= std_logic_vector(to_signed(-91,16));
ROM(4039) <= std_logic_vector(to_signed(-89,16));
ROM(4040) <= std_logic_vector(to_signed(-88,16));
ROM(4041) <= std_logic_vector(to_signed(-86,16));
ROM(4042) <= std_logic_vector(to_signed(-85,16));
ROM(4043) <= std_logic_vector(to_signed(-83,16));
ROM(4044) <= std_logic_vector(to_signed(-82,16));
ROM(4045) <= std_logic_vector(to_signed(-80,16));
ROM(4046) <= std_logic_vector(to_signed(-78,16));
ROM(4047) <= std_logic_vector(to_signed(-77,16));
ROM(4048) <= std_logic_vector(to_signed(-75,16));
ROM(4049) <= std_logic_vector(to_signed(-74,16));
ROM(4050) <= std_logic_vector(to_signed(-72,16));
ROM(4051) <= std_logic_vector(to_signed(-71,16));
ROM(4052) <= std_logic_vector(to_signed(-69,16));
ROM(4053) <= std_logic_vector(to_signed(-67,16));
ROM(4054) <= std_logic_vector(to_signed(-66,16));
ROM(4055) <= std_logic_vector(to_signed(-64,16));
ROM(4056) <= std_logic_vector(to_signed(-63,16));
ROM(4057) <= std_logic_vector(to_signed(-61,16));
ROM(4058) <= std_logic_vector(to_signed(-60,16));
ROM(4059) <= std_logic_vector(to_signed(-58,16));
ROM(4060) <= std_logic_vector(to_signed(-57,16));
ROM(4061) <= std_logic_vector(to_signed(-55,16));
ROM(4062) <= std_logic_vector(to_signed(-53,16));
ROM(4063) <= std_logic_vector(to_signed(-52,16));
ROM(4064) <= std_logic_vector(to_signed(-50,16));
ROM(4065) <= std_logic_vector(to_signed(-49,16));
ROM(4066) <= std_logic_vector(to_signed(-47,16));
ROM(4067) <= std_logic_vector(to_signed(-46,16));
ROM(4068) <= std_logic_vector(to_signed(-44,16));
ROM(4069) <= std_logic_vector(to_signed(-42,16));
ROM(4070) <= std_logic_vector(to_signed(-41,16));
ROM(4071) <= std_logic_vector(to_signed(-39,16));
ROM(4072) <= std_logic_vector(to_signed(-38,16));
ROM(4073) <= std_logic_vector(to_signed(-36,16));
ROM(4074) <= std_logic_vector(to_signed(-35,16));
ROM(4075) <= std_logic_vector(to_signed(-33,16));
ROM(4076) <= std_logic_vector(to_signed(-31,16));
ROM(4077) <= std_logic_vector(to_signed(-30,16));
ROM(4078) <= std_logic_vector(to_signed(-28,16));
ROM(4079) <= std_logic_vector(to_signed(-27,16));
ROM(4080) <= std_logic_vector(to_signed(-25,16));
ROM(4081) <= std_logic_vector(to_signed(-24,16));
ROM(4082) <= std_logic_vector(to_signed(-22,16));
ROM(4083) <= std_logic_vector(to_signed(-20,16));
ROM(4084) <= std_logic_vector(to_signed(-19,16));
ROM(4085) <= std_logic_vector(to_signed(-17,16));
ROM(4086) <= std_logic_vector(to_signed(-16,16));
ROM(4087) <= std_logic_vector(to_signed(-14,16));
ROM(4088) <= std_logic_vector(to_signed(-13,16));
ROM(4089) <= std_logic_vector(to_signed(-11,16));
ROM(4090) <= std_logic_vector(to_signed(-9,16));
ROM(4091) <= std_logic_vector(to_signed(-8,16));
ROM(4092) <= std_logic_vector(to_signed(-6,16));
ROM(4093) <= std_logic_vector(to_signed(-5,16));
ROM(4094) <= std_logic_vector(to_signed(-3,16));
ROM(4095) <= std_logic_vector(to_signed(-2,16));
                                                                              
process(clk)                                                                  
begin                                                                         
    if rising_edge(clk) then                                                  
        if rd_en='1' then                                                   
            for I in 0 to 8191 loop                                             
              if to_integer(unsigned(addr_in))=I then                         
                data_out <= ROM(I);                                           
              end if;                                                         
            end loop;                                                         
        end if;                                                               
        data_out_en <= rd_en;                                                 
    end if;                                                                   
end process;                                                                  
                                                                              
end rtl;                                                                      
